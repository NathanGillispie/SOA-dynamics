netcdf heatrestart {
dimensions:
	spatial = 3 ;
	atom = 3003 ;
	cell_spatial = 3 ;
	label = 5 ;
	cell_angular = 3 ;
variables:
	double time ;
		time:units = "picosecond" ;
	char spatial(spatial) ;
	double coordinates(atom, spatial) ;
		coordinates:units = "angstrom" ;
	double velocities(atom, spatial) ;
		velocities:units = "angstrom/picosecond" ;
		velocities:scale_factor = 20.455 ;
	char cell_spatial(cell_spatial) ;
	char cell_angular(cell_angular, label) ;
	double cell_lengths(cell_spatial) ;
		cell_lengths:units = "angstrom" ;
	double cell_angles(cell_angular) ;
		cell_angles:units = "degree" ;

// global attributes:
		:title = "default_name" ;
		:application = "AMBER" ;
		:program = "pmemd" ;
		:programVersion = "14.0" ;
		:Conventions = "AMBERRESTART" ;
		:ConventionVersion = "1.0" ;
data:

 time = 200.000000000591 ;

 spatial = "xyz" ;

 coordinates =
  7.32591327417033, 5.02903659894545, 75.1936341877445,
  7.364999297489, 6.00012157884252, 74.958121460701,
  6.89406864422518, 4.52220530663479, 74.4475562717583,
  27.3073357354856, 29.9783758312183, 86.2443679238097,
  26.6146145084018, 30.4535250519359, 86.7869271552296,
  28.173251689939, 30.4754344451006, 86.3002454164919,
  16.0559264909615, 24.9572587369228, 77.6425539504796,
  15.6076896673673, 25.8504514179682, 77.6066292444822,
  16.7365189941726, 24.8962337281894, 76.9124376632472,
  21.3471308923254, 2.77203061330173, 85.8470879675649,
  20.5182279901041, 3.29655864767654, 85.652690642882,
  22.0792887439997, 3.39533007965596, 86.1217562319755,
  13.0994396045212, 17.0738313101526, 61.3056919811106,
  13.5944817132361, 17.1438235617129, 60.4396467194062,
  13.0151099348334, 16.1116253271639, 61.5646285623639,
  24.7727822980166, 2.4332761085557, 90.00993113017,
  25.133294498856, 3.29529261556423, 89.6536187746577,
  23.8021032047381, 2.35814745826878, 89.7815941340917,
  6.50413032779126, 3.93719346333937, 57.6588074605006,
  6.22060177862739, 2.98370203412604, 57.5565056705566,
  7.48826023233912, 4.01145011720484, 57.4976420785747,
  16.2814196812407, 0.854505450512693, 81.3095842728863,
  16.3079186800068, 1.28595611061885, 80.4078370073188,
  17.1868488403026, 0.49369578402948, 81.533223317985,
  5.46110487338888, 28.7224674189762, 61.2831536564362,
  4.67999749459799, 28.838343319052, 61.8967040118106,
  5.59797947760828, 27.7493583008476, 61.0978863173427,
  30.941128056515, 19.3259116487612, 81.7755989975865,
  30.7984778288543, 18.3733785649425, 81.5066535816019,
  30.4940389290789, 19.9292723258019, 81.1152451488589,
  3.60945696787731, 21.7011995509675, 87.2864130002682,
  4.58104320083786, 21.4852590949143, 87.18951144527,
  3.0790194173675, 21.1455864809396, 86.646155144851,
  21.0152309090628, 19.5245493207828, 87.0981484835967,
  21.0796197399459, 19.1058494213137, 86.1923093849472,
  20.3036074172001, 20.2270723154082, 87.09083767983,
  15.6850096511919, 24.5158157365937, 69.8846634887508,
  15.3838618467111, 24.9431676330862, 69.0322080022762,
  15.910612442444, 23.5564718431205, 69.7150678678316,
  22.1839960277089, 17.0325179359001, 65.8379849865119,
  23.1762103885766, 16.9211779737197, 65.7821810896095,
  21.9681045819124, 17.7999480352268, 66.4416752434147,
  0.301893299615887, 22.960899825862, 68.3052263036995,
  -0.147949978283714, 23.85046445301, 68.2257542994744,
  1.25332699166556, 23.0921789760875, 68.5836858417814,
  25.6088697062717, 21.489823750051, 86.3866300214039,
  26.2394387862388, 21.9225390858514, 85.7423163760783,
  26.0446327899913, 20.6852778319355, 86.7901351645071,
  29.295376920623, -0.249292935921786, 67.1811805215803,
  29.6691259344832, 0.241454238862827, 66.3941107120466,
  28.9753685860722, 0.40858192169425, 67.8629395241133,
  18.5256882355682, 24.0889431056833, 61.7850047955393,
  18.189080152379, 23.3420112556521, 62.3584050133111,
  18.927183633986, 23.7131284539891, 60.9498013516879,
  6.8733008294904, 4.61431084052371, 70.9103289383499,
  5.90301352106751, 4.39722495931334, 71.0171758348541,
  7.4171257527069, 3.78625348246997, 71.0466207747219,
  28.0235322967807, 24.1858913915993, 88.5745459209939,
  28.6167259047698, 23.4446466194828, 88.2604161209895,
  27.0676099525501, 23.9358093802005, 88.420690601374,
  14.1348000102175, 27.0104332995846, 76.9893159258447,
  14.3598892683759, 26.999916670284, 76.015034536117,
  14.0721141664287, 27.9566347645799, 77.3067639887292,
  19.9846253635944, 26.0157868577294, 73.9072745330073,
  20.5631485881815, 25.2292309153641, 73.6913101189408,
  20.0251282944377, 26.6754388027715, 73.1567954700114,
  28.9227253970003, 0.9381982244869, 91.7655378164135,
  29.5432078321841, 0.78694895237853, 90.9960410943185,
  29.3868146218953, 0.702265361561047, 92.6193275302939,
  3.11593827014357, 24.2251128218139, 91.6427618075092,
  2.91367654395922, 25.1303711029036, 91.2691341336954,
  2.38675078759312, 23.5894095834911, 91.3894497310548,
  14.1937882481608, 22.432387585511, 84.9542524308183,
  15.1739673666805, 22.617951846472, 84.8848636660788,
  13.8013145459458, 22.9842535379111, 85.6900569997434,
  18.0301445376456, 11.610343104334, 85.2951773538293,
  17.8355524655854, 11.7505171518194, 86.2659941037378,
  19.0075694188572, 11.7407060210656, 85.1289061550914,
  23.0036997000513, 24.866903490204, 60.7620279129531,
  22.720279533248, 24.0035046996221, 61.1794192610557,
  23.1592647768499, 25.5478652634557, 61.477632950841,
  18.5243811895829, 13.4187920034036, 62.1956267026325,
  17.7054473680114, 13.6009849634542, 62.739826225964,
  19.171818247429, 12.8823492450496, 62.7369717156669,
  19.4236590430501, 24.6229492309527, 91.7843510710438,
  20.2808760112143, 25.130453874875, 91.6970693095543,
  19.6233671584105, 23.6551582501761, 91.9376393164727,
  21.7208670717539, 20.3600843761428, 60.294513649032,
  22.4580366137806, 19.6948336966834, 60.17609659035,
  21.0298047189749, 20.2216729040796, 59.5850948101413,
  6.28446227794541, 24.8439725817659, 82.2157692288716,
  7.17978866984034, 24.4077028832834, 82.1259950557346,
  5.72369873029708, 24.3245531789883, 82.8605542532378,
  21.8033655880759, 26.3089020513519, 90.8143732621625,
  22.119478903699, 27.2122823816874, 91.104159994862,
  21.2633285786127, 26.3973630687488, 89.9773937661107,
  27.4815927660154, 0.366875081846325, 75.9926858217126,
  27.4709941784982, -0.439078674999146, 75.4008022083482,
  26.5938130476419, 0.824969300116675, 75.9479995952893,
  11.36045128137, 22.9385082341809, 58.430033032603,
  10.3744358583025, 23.0015520395651, 58.5843024854309,
  11.5321458091036, 22.6021665137546, 57.5040766425678,
  9.04633580369107, 16.7540856534801, 71.4352930124748,
  8.86035800972126, 16.3078843914405, 70.5598978480465,
  8.86171249019875, 16.1143552653105, 72.1813890267836,
  11.0879442261342, 13.4705002067638, 66.8793610425716,
  11.6419202319261, 12.6746846212845, 66.6348449103529,
  10.3413484248665, 13.1850256495009, 67.4802761669319,
  29.9605943759342, 16.3071322535782, 78.9158239165916,
  30.9583645537145, 16.2864261115029, 78.8523737155461,
  29.6889965280349, 16.3770958775621, 79.8756883342754,
  1.70901092783333, -0.0312248729755495, 67.9232693122728,
  2.16397709198511, 0.766045709371561, 67.5265762218352,
  2.30212527597201, -0.443790027485459, 68.6146486316889,
  28.8959030519629, 26.944112745551, 61.4549165601707,
  28.8460707805214, 25.9785701977122, 61.7103462628991,
  29.3835540145946, 27.034467372138, 60.5865660663615,
  20.394960020341, 18.87480217346, 72.03265376551,
  20.822297095738, 18.014744035967, 72.3113705108327,
  19.6506240645846, 18.685053580967, 71.3923730016141,
  14.6249885386501, 22.9684708953987, 79.0041056360676,
  15.1590871305363, 23.383735788566, 78.2676996592804,
  14.823548166213, 23.4369668947643, 79.8649689079526,
  29.9862830049592, 15.2293532199257, 60.2673756293618,
  29.7159698098768, 14.2752260664418, 60.3961084983156,
  30.9663721905986, 15.2749830412289, 60.0741319810821,
  9.43043772657829, 13.2502907018026, 88.0265477651572,
  9.05454816440314, 12.4938989244326, 88.5618780521528,
  9.63805460388596, 12.9329429434616, 87.1012447701696,
  28.1524795570822, 8.51676161672397, 59.6541781578307,
  28.3498036010995, 7.54682267372005, 59.5117644348364,
  28.3364433039866, 9.02168712263764, 58.8108469220148,
  26.9946693115374, 20.1107476269462, 68.255779017529,
  27.5369804789942, 20.8034737431887, 67.7803538125524,
  27.4285980943075, 19.8891710732906, 69.1290542561301,
  18.9912681355654, 3.32506353772536, 84.5278848938066,
  19.1480226974394, 2.8370876611151, 83.6692187472874,
  18.9575684608355, 4.30870797748791, 84.350944372593,
  0.46553917864119, 29.840540490756, 64.0410628817708,
  0.0663390232104852, 28.9919206846787, 64.3881704452687,
  0.160723532961697, 30.6076315796552, 64.6055614942406,
  8.12625333732861, 4.09668119722868, 79.4066039063371,
  8.79856883670842, 4.72141669360025, 79.803715262089,
  7.22081534716624, 4.52029595582438, 79.4336701633862,
  8.49623444768988, 19.2427830395206, 74.6342734292674,
  7.87674262475782, 18.9092707126349, 75.3449065337141,
  8.99043345771429, 18.4711368442885, 74.2338617812416,
  8.4488977805755, 18.7219576715097, 89.5003755039138,
  7.53526426964094, 18.759638960612, 89.095586758827,
  8.93076894551776, 17.9140806121006, 89.1610602562787,
  15.1679359876969, 2.86457491946972, 83.1437473314324,
  14.5765913530074, 2.99549277169882, 83.9394684125856,
  15.1613798155359, 1.90039256682349, 82.8785881199156,
  2.91190147307633, 7.44516752754543, 80.1725532835806,
  2.00858174685209, 7.4601334737321, 79.7438465158839,
  3.52720693369116, 6.86996608475398, 79.6335333485613,
  19.3444464127563, 23.0215084450943, 85.0674841774561,
  20.1891628967732, 23.3302511595096, 85.5046706341605,
  19.5626460807946, 22.3573642904847, 84.3524307201777,
  29.4573504733679, 27.8811619710308, 84.6846072777431,
  30.0013206253057, 27.7610686416434, 83.8541411038158,
  28.5224132110409, 27.5673803428461, 84.5189769504287,
  14.6549701180719, 5.52005368517035, 80.9283567459752,
  15.5774484874289, 5.39779009668457, 81.2945333058462,
  14.6503874758548, 5.29429525209783, 79.9541842102881,
  22.5515013975177, 7.92162116086212, 60.8764757903549,
  23.3962447406834, 8.30012950305195, 60.4981371601968,
  21.8520577052883, 8.63551883624201, 60.9100708865414,
  9.94296549958411, 27.9288040183975, 59.492347315766,
  10.0711088258409, 28.7376501233531, 60.0662351675575,
  9.82095168024721, 28.2111326396693, 58.5408205544494,
  8.22423159454764, 27.9338661770703, 80.2237288273916,
  8.27716921121145, 28.0155147557498, 79.228474529063,
  8.4823610168524, 28.803887301436, 80.6437674500182,
  8.71293451811942, 29.0202291690905, 86.0234800370717,
  8.32698710934483, 29.9366464690358, 86.1294230879108,
  9.2120725893547, 28.7707590969877, 86.8533148814646,
  6.92412795907053, 7.6945688938615, 74.4180491694186,
  6.37153260611317, 8.06716910924735, 73.6725242165268,
  6.59571736252968, 8.05759587045936, 75.2900342004495,
  19.2380515254812, 13.7943921990013, 74.359723805456,
  19.5121153698493, 12.8384285645181, 74.2547355263205,
  19.471759453097, 14.1090569689349, 75.2797057004584,
  22.8352725145992, 10.891836280054, 89.2932762586413,
  22.1203277902313, 11.5186836385598, 88.9835724804389,
  23.7301757073113, 11.2476721854004, 89.023964015808,
  8.32681856071629, 7.44234217167192, 59.4370593984529,
  8.54338462908605, 6.60062483754784, 59.9316411080479,
  8.71699785137993, 7.39836447900354, 58.5173713623859,
  17.7013638525561, 22.8002947910477, 89.5752120683468,
  18.4925776810698, 22.7747461719045, 90.1862177521408,
  17.3550103296648, 23.7366097413479, 89.5173022157723,
  15.9382709428424, 13.3914484320251, 74.7069503978362,
  15.709905170215, 13.9959151857488, 75.4701469764023,
  16.3653859240293, 13.9239762205356, 73.9762062926189,
  26.5062337526509, 5.73709368755872, 74.3559087976037,
  26.3622812445953, 4.7507072456187, 74.2764137500761,
  26.0765154773088, 6.07010969550695, 75.1952195519059,
  29.7560903131012, 17.6020315948817, 71.5955291396928,
  30.3366627506626, 17.0619530888476, 70.9862255601333,
  29.0197608618882, 18.0242257595358, 71.0667843746044,
  19.7875873915216, 28.6020720078373, 86.0797936431916,
  20.0911891554193, 29.4664789536112, 86.4805761291564,
  20.2399271436836, 28.4662457809039, 85.1983516515149,
  25.1105424926282, 29.6347198639169, 83.9857074416172,
  25.8781884944834, 29.6132124891201, 84.6262205551949,
  24.6018957348964, 30.4875968282074, 84.103518135663,
  18.4240382140885, 19.6395665970204, 84.2542449665702,
  19.3611075587183, 19.4129864193949, 83.9886090005146,
  18.433578716784, 20.1258913484626, 85.1279710191421,
  21.792256634783, 15.098901788496, 60.9509968001638,
  21.241304649181, 15.5525116063617, 60.2505040859283,
  21.5679989573835, 15.4780263768455, 61.8487568129937,
  7.72141613598015, 1.98443221215858, 91.0282467655908,
  6.75373328904411, 2.10124431031236, 91.2517301910851,
  7.92984710028933, 1.0096369098595, 90.9486813727822,
  18.8429747687296, 16.3155428013739, 87.4438171327239,
  18.3609101230729, 15.4395248820856, 87.458179670586,
  18.9206939350921, 16.6685836381778, 88.3761914667382,
  6.41175398361524, 22.63022224966, 60.111442110759,
  5.48653682124859, 22.3474495223669, 60.3644495951571,
  7.03692665129513, 22.441038945978, 60.8686533185432,
  13.2626232214343, 16.343402551527, 73.6703855553443,
  12.8545980646192, 15.9928937680539, 74.5133915245487,
  12.8179269810659, 15.9172949972526, 72.8825546052081,
  24.9215751346551, 12.7862668435086, 64.0578446724842,
  25.6532829651291, 13.3286062294807, 63.6449625570488,
  24.1221046471696, 12.7929585984934, 63.4571765777305,
  25.1280995188614, 24.836035376604, 77.4603576921935,
  24.3591122134428, 24.6051142258509, 78.056456632169,
  24.7974641695139, 25.3676030547419, 76.6805397202789,
  6.71805990699908, 0.464948976826825, 66.7729906344426,
  7.19496273313445, 0.732585548207387, 67.6102088617189,
  5.85145468195873, 0.959980447767612, 66.7102273751982,
  28.9511179336606, 21.8523182036288, 67.2557457381836,
  28.3552764335261, 22.536858486598, 66.835772515573,
  29.7492369434156, 22.3044062535509, 67.6540200674911,
  9.68126664750307, 19.145667452022, 64.8968619199744,
  9.43608206755857, 18.1764970000053, 64.9212167284331,
  8.85854600554363, 19.6939830282728, 64.7469260198884,
  21.086393580738, 31.352617013303, 71.2894965224962,
  20.6475140352233, 30.4581398721708, 71.2040834759472,
  21.8831113271983, 31.2771162227919, 71.8891134528004,
  19.3009557385407, 14.0767623731042, 90.2601405242144,
  20.1394273826328, 13.7213869101382, 89.8470139305714,
  19.4160812534169, 15.0488734326591, 90.4644594017456,
  10.4412110789955, 27.7120166617136, 91.1225790865799,
  11.3191610213321, 27.5464558714371, 90.6733647463433,
  9.87283191931381, 26.8919452640923, 91.0560356147514,
  22.972811675267, 23.8311714716895, 91.340479825076,
  22.667614177477, 24.7714859943015, 91.1899371869044,
  23.9235325424971, 23.8348779500114, 91.6505057830725,
  5.5549261719187, 6.12393135382461, 64.1005446337865,
  4.89040378650283, 5.63697182439245, 63.5337286001597,
  6.42075927856476, 5.62360656563192, 64.1033973089494,
  28.8356031503367, 19.4498332267599, 89.0064077601108,
  29.3666040863155, 20.2617281613233, 88.763787436931,
  28.2639145086676, 19.6508662009992, 89.8018685324026,
  19.1016290391004, 23.3957408600349, 72.2556037021736,
  19.7988377888695, 22.8478560791389, 71.7933026897282,
  18.323592739509, 22.8139916887539, 72.4927269153604,
  10.9629541698489, 12.0806274380882, 76.783445123777,
  10.1327582159322, 11.5629107293499, 76.9901915568624,
  11.659125493784, 11.4624162394846, 76.4185336253947,
  20.896558717038, 11.1910573680874, 77.7083938974994,
  21.5343860139097, 10.6630598036221, 77.1476846044748,
  21.0065399946559, 12.1651420649824, 77.5107499705794,
  5.91605192218728, 30.2906194687761, 84.2192481741607,
  6.32352032304653, 29.5545885176702, 83.6786670596964,
  6.38563457202848, 30.3568626544072, 85.0996480692797,
  25.1878517532069, 0.41107124780816, 87.5063178894093,
  25.4569577707331, 1.30337292414213, 87.8687812251314,
  24.8009306911884, -0.144707530179929, 88.2421181623805,
  5.40519736499565, 13.5982618311324, 64.3268823610814,
  4.90710483228946, 12.9641454731857, 63.735443206606,
  4.81086009557001, 14.3652669059738, 64.5686806765001,
  29.8677585959786, 28.6219317488468, 87.373708518152,
  29.8132295228889, 27.8921006507021, 88.0551578180775,
  29.810259818256, 28.2268886787366, 86.4568470982425,
  19.7269939265003, 4.67968547655562, 79.8031799058567,
  20.0730361054467, 3.87347029077884, 80.2830464337714,
  20.2397549469642, 5.48703692356423, 80.0951726744416,
  23.3288248679889, 21.9386535944265, 64.7000934550052,
  24.004199674578, 21.7823871318362, 63.979364890777,
  23.7590676828235, 22.4256330389184, 65.4601869630195,
  25.5669999292079, 21.7140192773579, 76.5971610027624,
  26.4574274400171, 21.2655973273577, 76.6749851812179,
  25.0166372030918, 21.5048214573578, 77.4054537355078,
  8.14137815505856, 10.2637569405341, 82.8614399711104,
  9.04405176861021, 10.0299929971181, 83.2227359248051,
  7.98643398789699, 11.2465677443337, 82.9618154113212,
  3.38337037055626, -0.151675878611089, 85.1508103858517,
  3.57058089062856, 0.68963354460557, 85.6579106477143,
  4.11180386329662, -0.307916784744491, 84.4837471010693,
  8.91228359389411, 8.02920390696107, 67.8558474514086,
  9.16357336634285, 8.70480297320276, 68.5489703495703,
  9.38209046848626, 8.24041507443142, 66.9987177393336,
  18.0296144182193, 11.0041764945639, 69.0724976033063,
  17.6788094418998, 10.1776894575436, 68.6322078734388,
  17.4099565168117, 11.7675996200881, 68.890263642042,
  22.307715699965, 6.99012267970815, 74.2410525474414,
  23.0563325806166, 6.56967028184048, 74.7536855030059,
  22.0240962263533, 7.83377262737848, 74.6969195894439,
  25.6280639189496, 8.56768207530953, 85.2599551498717,
  26.2034094308133, 8.9802128170028, 85.9662100111904,
  25.0281470089958, 9.26569849276918, 84.8689656588258,
  3.17561308122482, 20.253098580488, 67.9293383651499,
  2.6750094142805, 21.0809520912804, 67.6762483943675,
  2.52863764223852, 19.5063205339284, 68.0834335647021,
  15.0925236786252, 21.0926979506602, 75.6390947348271,
  14.1101721138255, 21.1511669455767, 75.8167651594036,
  15.501629561041, 20.4134518587726, 76.2484034608668,
  15.4204488592156, 18.1974147540097, 72.4199588384156,
  15.248090019809, 17.2869117108602, 72.7958266860614,
  15.2506121998636, 18.8865009204685, 73.1244556548281,
  27.6498131445212, 25.085432716375, 78.2866028790457,
  26.7581250839626, 25.0456256633319, 77.8357062155126,
  27.9637044678201, 26.0342544518451, 78.3213814853591,
  28.7420633104747, 2.17847298606858, 79.0649240085301,
  29.598939504955, 2.62966673254906, 79.3142980057107,
  28.0756257627057, 2.86544309625638, 78.7752119745512,
  5.13860291322262, 6.16963345744521, 79.0193329378239,
  5.03683203817084, 6.05047198413367, 78.0316876410349,
  5.01316138216062, 5.28890233629148, 79.4760353732413,
  13.061581222052, 15.7735203799631, 82.8313971452946,
  13.9817145681374, 15.8880509518321, 83.2058799533501,
  12.4647015985317, 16.4922377459985, 83.1880202836149,
  1.67691810405885, 1.91850829989444, 82.7134160661332,
  1.40225626166943, 1.13674548472568, 83.2732444087122,
  0.99618230455173, 2.07099686987882, 81.9969343794912,
  16.2438487125763, 19.6593090736423, 65.8872009232909,
  15.674994513304, 20.0574889312807, 66.6068242281813,
  16.0102350828922, 18.693634416146, 65.7736354008144,
  23.28209625617, 5.08116641820667, 76.9483918821265,
  23.9557909436395, 5.42252575305128, 77.6038377399895,
  23.5024771409076, 4.1365386340605, 76.7052651352198,
  7.91753371362607, 7.43803009143006, 82.1172562280009,
  7.53817895245599, 7.69682928874087, 81.2289359362993,
  8.02029939130456, 8.25388359046461, 82.6863100774777,
  15.1034809445868, 23.0765244720311, 61.2670413043881,
  15.9013705052895, 23.3249852199545, 61.8162584797049,
  14.7953684212649, 22.1600624856314, 61.5223139046734,
  12.1408186998856, 29.1288125587596, 80.1321350131048,
  11.5015349349227, 29.5056004573089, 79.4618014040998,
  11.9550536627035, 28.1544277072703, 80.2588848144812,
  21.5511845167218, 3.76908561803926, 92.044125025641,
  21.7398956810467, 3.30186222028139, 91.1803597837802,
  20.5779428854409, 3.69035755824276, 92.2600014248659,
  11.7899098835425, 29.46083272939, 64.0322108284487,
  12.0596655661237, 28.5093909265316, 64.1805023234471,
  12.4027529673068, 30.0644321953382, 64.5422020434605,
  8.93786651683908, 30.4838567936167, 81.5511462989604,
  8.97990703369406, 29.9863084457217, 82.4175631942536,
  9.29068038671645, 31.4104416117052, 81.6813881820473,
  18.9422578534626, 6.71284487776283, 91.5513320156538,
  19.8880909490814, 6.94955070353643, 91.7735258663267,
  18.8991829204798, 6.35076302301547, 90.6201815011765,
  2.53517174992176, 27.1641329794016, 60.8158559506734,
  3.42040034123538, 27.2851502581858, 60.3667177098649,
  2.56024750650246, 27.5874021069169, 61.721512868123,
  12.4889817624226, 27.6534914402749, 66.4008822858449,
  13.0795272187329, 26.8466589843839, 66.417539180878,
  12.191702707294, 27.8682621482857, 67.3312041153009,
  26.6387005031898, 0.216502365546534, 90.3510356550827,
  27.4124772339081, 0.42370633765071, 90.9496474532818,
  25.8922217618234, 0.855092743053374, 90.5380431908764,
  22.3578379687356, 1.65810613806948, 67.5847371078105,
  23.1842074910105, 1.53394384596142, 68.1340067482182,
  21.5517913904409, 1.49494922463394, 68.1536560257747,
  2.14201260967124, 15.0152417442114, 85.351476322771,
  1.37461598581043, 15.0180000928795, 84.7103095634956,
  2.99802979599475, 14.9052758100145, 84.8463604251445,
  28.2021810357388, 3.96341267352643, 70.9438509316534,
  28.3744423072986, 3.25006996059934, 71.6231654598614,
  28.3317724734101, 4.8617467075162, 71.3636151781751,
  24.2444187942858, 15.4148723799483, 76.2196900726618,
  23.7012810407271, 14.8048305493143, 76.7966219105212,
  24.0402409419748, 15.2333415106558, 75.2577347992111,
  24.0456275687684, 13.1795704174808, 84.5057569936043,
  24.7965830271692, 12.5281433369477, 84.3975504399847,
  23.1941278642723, 12.6821380555758, 84.6716162670039,
  21.0639486487685, 11.3582397877954, 56.2315427302735,
  22.0312115749534, 11.4084669351601, 56.480298966971,
  20.6189956536359, 10.6401311630275, 56.7666472389039,
  31.0014661179521, 0.968778606417392, 69.9165986799949,
  31.5709791311372, 0.527852644988917, 69.2228846003113,
  30.2278641559108, 1.42213333469851, 69.4738690845634,
  21.5493482651099, 28.8089014742297, 62.9423085307299,
  22.146647072227, 28.0099343653819, 62.8724107911669,
  20.5954389128302, 28.5201339538235, 62.8606368294392,
  20.9151297013134, 7.13918212815653, 63.0789603827782,
  21.1127382288239, 6.24340419156122, 63.4771221064084,
  21.4569453128789, 7.26120278301005, 62.2473674518,
  22.0981612678422, 13.3601770637034, 76.2975808005728,
  22.9739136241637, 12.8774248235645, 76.3004242207518,
  22.1323370361907, 14.108783192527, 75.635447218321,
  26.3352532609847, 20.6292479469757, 72.027940664694,
  25.9047642410553, 19.7298250933681, 72.1035563649732,
  25.6430117655536, 21.3113920753023, 71.7923964009285,
  21.6522421801735, 17.1575066683404, 82.0273634955123,
  21.7621399415644, 16.4996965989887, 82.7724865690383,
  22.4710240399979, 17.1507834970197, 81.4532981116143,
  3.39176063424484, 20.2868978052909, 74.6801763884516,
  4.27922285215538, 20.7355595853338, 74.7855965900736,
  3.27205337112967, 20.0043350042883, 73.7284261929449,
  19.8150510715182, 11.2646786750032, 63.0611768374088,
  19.1386724783287, 10.5603328080265, 62.8457495913422,
  20.545326449289, 10.8668151911137, 63.6165168420988,
  0.14752269599001, 18.8301161155683, 73.2917033482449,
  0.967870345658872, 19.0517305850863, 72.7645252373725,
  -0.46310651645317, 18.265469821293, 72.7364497779977,
  6.96924406879072, 6.53606554315825, 56.1706089989926,
  6.16390824942135, 7.03145527283238, 56.4962210899444,
  6.87021869376318, 5.56358229803414, 56.381488853539,
  27.4616587759319, 30.3235493751108, 62.2493418644388,
  26.4821508945453, 30.2227696592622, 62.0749636571563,
  27.9554094055983, 29.5635460115485, 61.8267247764288,
  27.5901004926904, 4.68029667727253, 85.3555861918686,
  28.3271479964821, 5.34813086278308, 85.4593092742459,
  27.9732444636469, 3.80336839548036, 85.0654181610438,
  22.192826886023, 10.7731607571863, 71.1837338867187,
  21.4477972847955, 10.6889330772129, 70.522041668825,
  22.7769367922094, 9.96307641688515, 71.1329502368524,
  9.49600059753297, 4.30701975313439, 57.7516797681097,
  9.85396787381596, 5.10768921989088, 57.2712759441091,
  10.2482851736402, 3.82168736333794, 58.1972360361226,
  21.492024790428, 15.9509069190972, 78.9382474554185,
  22.056688074641, 16.7617870535623, 78.7845308883495,
  20.5661431117302, 16.1205692417461, 78.6006710739502,
  19.77750946473, 14.0374707056862, 84.0131868978463,
  20.5923783892076, 13.6252353732352, 84.4206800469908,
  19.5459301400588, 14.8759449726705, 84.5064737515024,
  18.64292481407, 30.9730817364067, 82.4070957932734,
  18.4232007399715, 31.1805182221286, 83.3603488738627,
  19.455807722434, 30.3917571958701, 82.371274628305,
  26.9319656739396, 28.3754497956018, 67.6218892703721,
  26.8853711784191, 28.2313246658582, 68.6103511563159,
  27.195396351864, 29.3218647469713, 67.4350657767947,
  25.8549652591388, 8.55556547251056, 90.644488770165,
  25.8362583331879, 7.60479168024338, 90.9538093916234,
  24.9928699277527, 9.00146107538233, 90.8852557756744,
  26.53648015176, 3.6807808199478, 61.5721483390119,
  26.0472828026302, 4.55232231083575, 61.6053354338714,
  25.9388556434754, 2.97751888180279, 61.1870930268111,
  24.1400628759739, 22.3143605527471, 71.3028588357542,
  23.621681705393, 23.1111232306334, 70.9922945153396,
  23.8987002262945, 22.1086137457808, 72.2512323501265,
  2.44772493982272, 19.4969278001756, 85.8593926669006,
  1.76182524126784, 20.0744540244601, 85.4166680755507,
  3.21280271685683, 19.3481083395984, 85.232887468804,
  8.85096685396785, 24.4931330358976, 90.5386918814207,
  8.84402426123124, 23.5641208042049, 90.9086757645447,
  8.01116246214865, 24.6514093287062, 90.0193873478222,
  14.1272074308216, 30.1269884860192, 65.1919337324511,
  14.4318339491637, 29.1761920047183, 65.1354648430651,
  13.8463430789779, 30.3319110902336, 66.1295487612051,
  17.4416968082606, 9.2970198998268, 80.8363794166318,
  17.077575959692, 8.75849709991626, 80.0765049522535,
  17.2730926922364, 10.2681490497729, 80.6676167839649,
  13.7179654357851, 29.5744039706148, 91.3438466734157,
  12.9956046489736, 30.1927511602098, 91.6534296942632,
  13.3068136218769, 28.756147617273, 90.9420871357121,
  1.80318618841121, 11.3338891661268, 71.7659456191607,
  2.65542831116705, 11.0737220075377, 72.2198138971801,
  1.02588299239037, 11.0150505601512, 72.3082939249526,
  8.99520688019007, 2.44126661051132, 81.6653409154681,
  8.45847215628121, 2.77306849806625, 80.8895681758301,
  9.54220425669643, 3.19120861407303, 82.037336696881,
  26.225547836083, 24.4440908399253, 71.4524220473093,
  26.9804043250236, 24.138197221638, 72.0326123397095,
  25.5136524942073, 23.7420481877234, 71.4339521608722,
  17.6267236802812, 21.6857575650745, 62.8801040292561,
  18.4387613728203, 21.1184415934589, 63.0170250803975,
  16.8135413031621, 21.1780529508905, 63.1646570933393,
  3.09543873820108, 23.0826574847779, 68.7954978706842,
  3.20468330175341, 24.0737776268878, 68.7196922690558,
  3.28725472987991, 22.7969983137727, 69.7344363475595,
  23.7106301290555, 18.1617928412959, 76.962780319331,
  24.1863472143198, 18.4489603313674, 77.7941815987585,
  24.1363791027336, 17.3305422090548, 76.6053447337904,
  12.6947306544931, 13.491139614298, 87.8802814204996,
  11.7355951070901, 13.2745664499935, 88.0623667472316,
  13.0381722537246, 12.8974692917853, 87.1525428574943,
  16.1703647792341, 13.9108059288646, 63.3942070849497,
  15.4336612003733, 14.5853565348461, 63.4416340484169,
  16.4163129746984, 13.6202281764379, 64.3189092288547,
  8.72570417486004, 2.19470121324143, 77.4265905527985,
  8.45250309790054, 2.90517265218998, 78.0751208188512,
  8.07514649234018, 1.43644154636044, 77.4692165929139,
  30.5786738733154, 23.576788239276, 91.0080726677933,
  29.8461010752481, 23.4113442119575, 91.6683494047427,
  30.9744277563274, 24.4809599287041, 91.1688595457332,
  19.6342029704358, 22.7750031766188, 59.3668288644391,
  19.8625292992556, 22.018041418207, 58.7545576958627,
  20.4700908114956, 23.2607518973859, 59.6224451734679,
  29.7056029167102, 19.7631361122814, 65.4075332717706,
  29.8775000585269, 19.0959327552111, 66.1323029268676,
  29.2435017415539, 20.5619968190653, 65.7926099850056,
  27.3862560378392, 9.75309978801125, 87.3497302147071,
  27.8263183545567, 9.78891337881847, 88.2469829907511,
  27.9930032677145, 10.1560656068386, 86.6645467736524,
  8.36807486146038, 12.658096465829, 61.6869903670616,
  7.70010004382219, 12.5894621675399, 62.4280024965842,
  8.61905601374701, 11.7406092992462, 61.3784036525827,
  8.70141529617887, 4.87509120933911, 60.5055169537221,
  8.84942422056298, 4.51563248884033, 59.5841686012733,
  7.84416339580218, 4.51248119666481, 60.8710756466961,
  2.84811557955566, 19.1916877745674, 81.6763086417174,
  1.97801365100041, 19.671211443173, 81.7902370629806,
  2.67351772628514, 18.2309130189857, 81.4608383220205,
  25.8180480965285, 0.556176507887081, 68.3552763562186,
  26.1433542105932, 0.771581413612978, 67.4345284761009,
  25.1150626039944, -0.153104596671792, 68.3030105738911,
  24.8957636924172, 16.9398685903097, 65.7651617210957,
  25.5634027991511, 16.3289282691482, 66.1906143590457,
  25.3655944211291, 17.7414953631439, 65.3954948393852,
  12.7721445870424, 5.68140994219371, 69.4365692786507,
  12.2432257991944, 6.31502614667195, 70.0011712812011,
  13.7484224189621, 5.85523898444704, 69.5656624967973,
  17.8055242189367, 5.39687480570711, 89.164615941025,
  18.0006027803923, 5.81586418248508, 88.277828335672,
  18.3456299670267, 4.56122650074249, 89.264504335195,
  4.59694044554109, 12.2851699392962, 69.271040589544,
  3.59865917607531, 12.2463312151305, 69.31492749578,
  4.91322435811949, 11.810379560188, 68.449737611009,
  2.65860442794997, 12.8754292594288, 79.5843058939994,
  1.7047189106103, 12.8836507181312, 79.2842478539031,
  2.92204426276563, 11.9431533169578, 79.8322192266826,
  18.0754530310693, 25.5047146126694, 70.7127654310052,
  18.3565970727734, 24.9241351675503, 71.4768894626384,
  17.1549078118758, 25.2468748751851, 70.4193115688835,
  8.59940715159373, 10.8871708826383, 76.0627218991936,
  7.95023150936911, 11.6012585708718, 76.3247328895271,
  8.93279345262648, 11.0632773323172, 75.1365253257465,
  28.0754862526183, 30.4192253028866, 82.7633052145145,
  27.9842366189807, 31.4135430372333, 82.8181299126404,
  28.3223933921529, 30.0570754105709, 83.6621290681936,
  1.06126219005576, 16.9067579996972, 63.634935191173,
  0.0950410037770014, 16.9931503258456, 63.8777375494167,
  1.33882259110982, 17.695212314478, 63.086027168577,
  15.0907225294755, 22.5186834792033, 88.201828956377,
  16.0237782748787, 22.3541582786864, 88.5217327456088,
  14.5666761347468, 21.6684142235879, 88.2509977384155,
  17.759297015017, 11.8014961663431, 58.1524128276947,
  18.3667214670135, 12.4904642286059, 58.5478348102635,
  18.3016889488013, 11.1266976243049, 57.6519551193629,
  2.79551156588106, 5.67272655159616, 73.5099406642669,
  1.80103423467985, 5.57917076831963, 73.5575027620174,
  3.16677032244209, 5.75937211209763, 74.4344186156114,
  11.2591105997637, 14.7933515160094, 64.4035429083646,
  10.6419131614356, 15.5696398012744, 64.5317763684349,
  11.1199084938037, 14.1315801971598, 65.1402120981943,
  9.73897676503542, 5.29808570366834, 82.3497240432627,
  9.25542758264468, 6.12912970508275, 82.624580471098,
  10.7092378335014, 5.3870716573573, 82.5748350360316,
  20.7317478116509, 28.8262862585054, 69.2734584943954,
  20.8682697632358, 29.5260643360007, 68.572264941236,
  19.9640044877292, 28.2402005312619, 69.0144725702697,
  17.2171336375206, 4.92523782901768, 79.0924662548517,
  18.1503875874783, 5.09263707656395, 79.4102941277787,
  16.9275109419597, 5.67593520878761, 78.4986884022649,
  26.7831816496143, 1.93105639827145, 65.9159381430043,
  26.3350374082986, 2.77696852113131, 66.2050737848306,
  27.7273080947997, 2.12759769653328, 65.6513691093305,
  8.34907022696572, 11.0489668318115, 58.3664522553196,
  8.6894159298248, 10.5267785618684, 59.1484268158259,
  8.73656151770416, 11.9706117740694, 58.3869729768517,
  31.2720556166317, 19.8551904902677, 69.6507089574943,
  30.3565350901286, 19.9023972112365, 70.0502007484575,
  31.5417616249097, 20.7621645261909, 69.3272019757151,
  5.43926503372422, 11.8703438111401, 60.2602563799514,
  5.52410067967822, 10.8764642193942, 60.3310113818006,
  6.23338398436826, 12.2391345691472, 59.7771741208727,
  20.9138987137102, 21.4089801821084, 71.1533886872673,
  21.5095847921847, 21.4128268772236, 70.3501805580453,
  21.0047307831082, 20.5354372524607, 71.6315855977879,
  20.2541070601479, 13.5178097090102, 65.5183333813466,
  19.2659731856064, 13.4407426459702, 65.6511946389728,
  20.7161003971084, 12.7877438520993, 66.0218867560519,
  2.35669387195217, 19.7327883751088, 71.627675476378,
  1.60515000136189, 19.6015149352815, 70.9811856508014,
  3.22604140601689, 19.7288073416815, 71.1334902718358,
  9.9289840849324, 3.63922379831085, 74.9407988606702,
  9.97899631449095, 2.68709554607997, 75.2423789797071,
  9.16005706129616, 4.09193249844548, 75.3922477117534,
  22.7668038996029, 4.16792996837353, 71.4466783148748,
  22.6371173645095, 5.15538839281963, 71.3566379761045,
  22.1176349664183, 3.69105848626158, 70.8540795587706,
  29.3460321689366, 17.0613444945019, 64.5428735801668,
  29.0155892276631, 17.3720639741279, 63.6516604364444,
  29.5538554724355, 17.8538956978034, 65.1161728603584,
  30.339546862753, 26.3917515414857, 91.61550481755,
  30.9611677015267, 27.1573500008614, 91.7811747659529,
  29.7406140947601, 26.6094093449913, 90.8448527430071,
  25.5182264056032, 17.5078911942955, 72.4590478138157,
  26.0155492054149, 16.656003643008, 72.2948600166171,
  25.5878696178545, 17.7535015931552, 73.4259114830883,
  12.6877008302198, 24.2130816091044, 86.454221143821,
  13.2550730676444, 25.0145225305821, 86.2650619685723,
  11.7691213609978, 24.5092271384859, 86.7159644993263,
  10.5483478595185, 25.9578873117721, 88.7025254618543,
  9.98970392305488, 25.9977909412243, 87.874078328593,
  10.1932691872708, 25.2474282175615, 89.3101166171292,
  10.5453556445871, 30.4543841171945, 78.2894025718898,
  11.0253175455564, 31.1648961812643, 77.7748064385685,
  9.66014433394912, 30.8047944192347, 78.5953658960687,
  22.6560232805059, 14.3734668265317, 71.2965829206482,
  21.7909938160427, 13.9687589609761, 71.0000435991949,
  23.1209932243811, 14.7796839217767, 70.5099504633828,
  15.3966688851921, 30.7942260271152, 86.9250066865101,
  15.4362518276575, 30.863085195073, 85.9281658739156,
  14.7962795279051, 31.5083760944405, 87.284898755047,
  5.07426836543336, 1.28151743702042, 69.579956750815,
  5.6781016183185, 1.03871282886326, 70.3391874963514,
  5.12869205138308, 0.577038209167302, 68.872321901524,
  24.4906408358354, 6.00075826525044, 88.8753032494841,
  24.711595595647, 5.65228941455273, 89.7862085432496,
  23.8118017637674, 6.73088786093629, 88.9533307301399,
  29.6138079392004, 10.7243705005491, 89.0794413104533,
  29.6440688962478, 10.1818182318501, 89.9189181178805,
  30.391305496906, 10.4833657424635, 88.4985676113224,
  24.8475664438615, 27.028978878936, 82.5808591227537,
  25.4422576450094, 27.1449861432864, 81.7853186210222,
  24.7630662272829, 27.9005439202305, 83.0638022790273,
  9.80794827637434, 11.7933343082425, 85.77037063794,
  10.3990793981387, 12.31238626443, 85.1529979274486,
  10.1605140244795, 10.8623627536399, 85.8651828617506,
  23.6480322780245, 16.0719440607953, 57.6570266668782,
  23.9114062150961, 15.3961122488936, 58.3454201090993,
  23.6254488453655, 15.6386588874352, 56.7560527787352,
  20.6971357908877, 0.293557955169944, 63.1083503549908,
  21.1737369946201, 0.679628790884452, 63.8981608401146,
  20.986453917661, -0.654349528214197, 62.9750596033808,
  16.3885947505324, 26.160105270279, 84.3015923472709,
  16.4378759272374, 26.6449402618277, 85.17480846977,
  15.667354133157, 26.5619932422374, 83.7374132712292,
  27.8568418412655, 24.3793751610046, 61.8879904092594,
  27.5303129685681, 24.4060540906873, 62.8328010410825,
  27.1319557271293, 24.029599363521, 61.2945285208224,
  1.29164634907628, 14.2468179445335, 82.6957596301379,
  2.00560555008037, 13.602913135652, 82.970803001992,
  0.656741195786527, 13.7933453071472, 82.0702534243589,
  29.2569882404139, 8.44394072613023, 69.2121432443698,
  29.6912897653217, 8.26279223413004, 70.0945079134884,
  29.7255262559209, 9.20261300507442, 68.7594971340514,
  7.24620658765911, 27.7693824639861, 93.3194174691957,
  8.0504318455319, 28.2651154923536, 93.6472444040028,
  6.42690359376476, 28.1328812798548, 93.7628261013374,
  15.9439607676454, 2.84033445400424, 91.0700867922597,
  15.0118894217265, 2.50013364564581, 91.1946115532886,
  16.496521373405, 2.14056464943084, 90.6173186423531,
  27.9880167832736, 22.3877629678378, 84.9345241314076,
  28.8536251082904, 22.6178680527342, 85.3792418818589,
  27.8462691526061, 22.9902806174063, 84.1491069867267,
  29.83587466511, 12.879357977728, 56.3394451328065,
  29.3805091448641, 13.6329893606842, 56.8134514424635,
  29.1504750404929, 12.2294328554218, 56.0110784323481,
  10.8145333815785, 23.7228899148515, 63.4278322943538,
  11.757712651097, 24.022791437682, 63.2847520995175,
  10.7125959910326, 22.7802770083167, 63.1098862661624,
  10.3813596297313, 16.0557096067691, 59.9495997417755,
  11.1796578729698, 16.391888442247, 60.449303359352,
  10.342396336374, 16.4925230144715, 59.0508918311492,
  14.8455593824768, 26.9368274691864, 71.5474282645805,
  14.8443103091764, 26.075451018257, 71.0394626657451,
  14.8947270301959, 27.7021823592747, 70.9057005694981,
  22.1207082802453, 4.68334689589041, 63.6694309307721,
  22.2016578649591, 4.88552005897768, 64.6454294844912,
  22.195529310332, 3.69650402640437, 63.5261027604728,
  7.07930658804272, 22.4463671950018, 89.333868003908,
  6.81329928906212, 21.6648633647786, 88.7695171553789,
  6.62112673147145, 22.3883566379054, 90.2208324870175,
  1.7876484366175, 10.9158744163375, 68.9738895175148,
  1.01947622897255, 10.8784013602492, 68.3347438146666,
  1.44021827262001, 10.9901640760884, 69.9086479502656,
  25.7929560052829, 23.1398218574017, 80.7537192813704,
  26.0931494276211, 22.1995044120986, 80.5934476018902,
  26.1366449509984, 23.7287232863681, 80.0222324287515,
  9.7190058569889, 25.2521966655775, 77.4206369267004,
  10.0386204728158, 25.3273510966481, 76.4760744307054,
  10.5049912515908, 25.1628711656976, 78.0323949789921,
  5.19064202080502, 26.0809307487452, 60.2675385956705,
  5.85726871294461, 26.1127101538518, 59.522824608466,
  5.10029248485806, 25.1400927075685, 60.5941281570913,
  24.4289292864283, 2.27662342631242, 76.4507337079773,
  23.5838135226777, 2.10544438952583, 75.9442980425419,
  24.2971762438297, 2.03223554563015, 77.411418723756,
  1.92576013492167, 29.9043002073952, 73.326854159821,
  1.17970458389374, 29.8375246501334, 73.9893812458581,
  1.78089153897234, 30.7016203544638, 72.740941476065,
  21.302687783061, 4.33887120287287, 67.2254702038596,
  21.2244184454524, 4.78312865107674, 68.1179438620175,
  22.0363242207114, 3.65993930541393, 67.2542635358027,
  27.5037533121935, 10.6487851903455, 91.5026663091242,
  26.9891906457687, 11.5031898611855, 91.5749014859327,
  26.912085865438, 9.93379561140092, 91.1302155950015,
  6.52384341384963, 14.6807772710447, 87.4270234054947,
  5.52903490812246, 14.5954869332695, 87.4825355232264,
  6.94697726159038, 14.1137553531392, 88.133736849198,
  27.5514956498243, 12.8145988585161, 68.503763312824,
  27.9357975317287, 13.6927671833501, 68.7886009101018,
  27.9660106608745, 12.5344509036577, 67.6379143485106,
  11.0420876607303, 6.04656287549469, 62.1549916127353,
  11.7255829409755, 5.48172551343032, 61.6926141086342,
  10.1288304431664, 5.68453501538339, 61.9681840029584,
  14.8150437911486, 12.2620117622518, 77.9205053081029,
  14.2837733079776, 11.6944148707424, 78.5494611431662,
  14.2256895055424, 12.9702424222664, 77.53182696004,
  21.5449640437627, 2.38624583701911, 89.55655949507,
  21.3167545149456, 1.42454607962447, 89.7083948914179,
  20.7675865050689, 2.85028736861522, 89.131883595956,
  2.68650647203482, 10.5037224203137, 86.0620794618555,
  3.49357676855831, 9.92092287082862, 85.9673048788208,
  2.71199064945771, 11.2237563133661, 85.3686086625013,
  29.5521501895229, 0.567703511509323, 86.241757163223,
  30.2066262674971, -0.109350748364428, 85.9052180235286,
  29.5546210186455, 1.36346295884783, 85.6361493718472,
  12.3411146442747, 26.426849498165, 81.0321464814747,
  12.3169623341489, 25.8578804321587, 80.2101423039649,
  11.4817814775971, 26.3251131494695, 81.5333412779381,
  24.1918149001127, 3.50074357848331, 93.1707140579208,
  23.2491457033281, 3.80866661624979, 93.0420354340306,
  24.3782669635253, 2.73287259366891, 92.5578439422116,
  26.79610572424, 28.3169339178627, 80.687027026671,
  27.4174301065084, 28.9078431460421, 81.2015970375065,
  27.2698010189764, 27.953172240131, 79.8849732818643,
  19.6986007125604, 27.4395392693143, 71.58059622903,
  19.9761557074466, 27.955178836178, 70.7699920951284,
  19.2765522747037, 26.5777679068152, 71.2991264528923,
  0.754824244851074, 24.73240435516, 63.7600569958326,
  1.6562724163486, 24.7394481496314, 64.1928867303278,
  0.338213089921831, 25.6377118676211, 63.8428425831652,
  5.69349465402708, 27.7060622046084, 74.7264619038579,
  5.86309546888485, 26.78221127008, 74.3833365413873,
  4.73212572201859, 27.7934481997859, 74.9874857809568,
  18.4174483726206, 21.1090851770437, 86.8729473175384,
  18.608427259472, 21.8825130310514, 86.2685166602898,
  17.9426038967625, 21.4343982606517, 87.6906845133297,
  27.8577559132831, 14.7738053026611, 57.8932411255127,
  28.4449417187797, 15.4243668400464, 57.4115954923984,
  28.1501469269186, 14.7035915464622, 58.846958863413,
  29.9770641238754, 1.06637711413499, 64.9065399885219,
  30.3089928673881, 1.74307130682595, 65.5637372791496,
  29.4649690828978, 1.52826362032846, 64.1823718282148,
  27.1204671734135, 15.1641012787423, 76.0671242997674,
  27.5636821383349, 15.7554508702047, 75.3934284072855,
  26.1294744351455, 15.2894473727688, 76.01998886286,
  1.46803923870723, 1.87521947915297, 71.9892158444699,
  2.0558504262516, 2.63122692551684, 71.7012388508748,
  0.968941872271668, 1.52108915921012, 71.1983343518844,
  11.4846519183818, 2.15903052955576, 63.8847375470774,
  10.8752285934694, 2.08122808966908, 64.6737559191071,
  11.911200609714, 3.06348699464241, 63.8809013137987,
  3.87458477552921, 2.02106868194975, 86.577942194488,
  3.54016834474175, 2.03437973352047, 87.5202735941163,
  4.75339170150197, 2.49576716386493, 86.5293650586139,
  1.5830510153638, 2.32107884652846, 74.6608711946074,
  0.904444171945964, 2.49333314551994, 75.3748888474321,
  1.1795460118306, 2.50852324300182, 73.7652996953096,
  20.3219220712805, 25.3186445186557, 76.5769563200023,
  20.3261479305647, 25.6851594501791, 75.6465537474114,
  19.5256698230925, 25.6694593511093, 77.0698166557832,
  17.4378980362998, 25.2107170045619, 74.9049684164966,
  17.0387251950847, 24.3406384553545, 74.6157896464503,
  18.3234883146314, 25.3361793047689, 74.4577670411059,
  21.4657547074293, 20.0753860801975, 64.8710220611431,
  21.3576536729513, 19.7683429035315, 65.8165582339084,
  22.096800816723, 20.8506016418091, 64.8423577805745,
  3.2280788138727, 28.8926166628926, 63.1343094348399,
  3.67796509533141, 28.3005006427766, 63.8028907331704,
  2.3300578732576, 29.1641457985473, 63.4804745958648,
  8.61307048074504, 18.7264332065378, 85.7787893029557,
  9.5248783114792, 19.0414953074473, 86.0421186639894,
  8.49805019509007, 17.7717763713495, 86.0533811107649,
  3.67209744206774, 4.38793021467182, 90.9587994508793,
  4.65418108383846, 4.31093081867445, 91.1307960019564,
  3.49642913094268, 5.18453238935193, 90.3803829748334,
  17.3931534766977, 13.9200211949894, 65.9060743789238,
  16.6997814290706, 13.5530638947595, 66.5262175425379,
  17.4401855376725, 14.9135917714913, 66.009057361742,
  31.0921286451106, 11.977494722413, 78.7557405462162,
  30.2627385358466, 12.3782894160831, 78.3665418049786,
  31.2462905596177, 11.0747713596626, 78.3540881660911,
  7.57012823142865, 28.3010886105676, 83.349522718267,
  8.03516494265285, 27.4636596473705, 83.0623753888134,
  7.95388875785346, 28.6143984380479, 84.218179618523,
  22.6789529277097, 27.0832870957639, 70.0535469283906,
  23.0803641507577, 27.4126682993566, 70.9081679278582,
  22.0119764496557, 27.749533668724, 69.7199935117665,
  3.74662454340026, 10.4137605827248, 77.8308515826405,
  3.4697618861007, 9.94012988085203, 78.6669263563519,
  4.28073985965858, 11.2250507042481, 78.0686102158317,
  26.9412078160497, 26.6234864981879, 84.2809405350001,
  27.1795729491016, 25.6656167094853, 84.1207296388788,
  26.0365502284204, 26.8104204278974, 83.8979909886259,
  7.19266487705974, 12.9326578413386, 83.0074273223537,
  7.6090264810371, 13.5346012463547, 83.6888281969429,
  7.31936755641657, 13.3233508687444, 82.0956678204123,
  12.244810281528, 14.4165456391497, 61.9256918978249,
  12.2018455797031, 13.6454976624483, 61.2903659562627,
  11.7966560734656, 14.1666176564113, 62.784000588938,
  0.327932322158198, 5.02849206202012, 60.0250408738034,
  0.900460153041788, 4.73817149937856, 59.2582776419181,
  0.420627911091259, 4.3751225233571, 60.7763835211619,
  14.1210803795536, 8.63963569658531, 84.7401145798307,
  14.9969613582588, 8.56544918671079, 85.2169047568426,
  14.2644409990802, 8.51536617797721, 83.7582771088032,
  9.57450231641331, 2.07668695047302, 66.1541945624116,
  9.49189222215113, 3.03309283890795, 66.4343076625925,
  8.67155447307887, 1.72063899298265, 65.9135391153828,
  17.1630540277821, 4.46593248159942, 82.0778722247956,
  16.4525019948658, 3.90310707389384, 82.5001794221763,
  17.4155877172008, 4.07519970341384, 81.1926860117534,
  0.444614260778938, 4.80479048548263, 83.396188338591,
  1.23216379105313, 4.20917918643184, 83.5543430660193,
  0.449626733087286, 5.54857025261439, 84.0645943029022,
  9.80412711962006, 10.2328968632421, 69.492269066216,
  9.55594883322871, 11.1197880874658, 69.1026134560179,
  10.7413119542342, 10.2716048939203, 69.8389479870207,
  4.12801793892036, 14.928597191367, 78.5072973068206,
  4.99517080655629, 15.1796246557937, 78.9374497405627,
  3.75655675795204, 14.1155790398443, 78.9556477014097,
  30.4902639784539, 23.1172055313973, 85.7570095443845,
  30.5022116187909, 23.4497325155725, 84.8139914858694,
  31.2192728854473, 23.5626004204541, 86.2767877724071,
  26.9013285404171, 12.2973161915803, 74.7507906723125,
  27.8351578364748, 12.190175128677, 75.0920876668266,
  26.7437276087668, 13.2538949180895, 74.5055987345717,
  22.1402789009978, 28.6102626229109, 66.0021963580411,
  21.9702358638946, 28.3799891967707, 65.044042135201,
  21.5746264579584, 29.3927704229888, 66.2624248278535,
  30.5889023283353, 9.71744262214364, 57.8669438943584,
  30.9578462505328, 9.12609846974189, 58.58401604951,
  31.2609872670333, 10.421188569968, 57.6366322010034,
  17.915906761377, 20.1139648784189, 73.5608545467088,
  18.0809718131427, 19.6853398098177, 72.6725786440455,
  18.7703718247047, 20.1461786909825, 74.0793636843645,
  16.9579196675117, 21.3036725446971, 82.2859039306613,
  16.7512242259272, 22.0051654141487, 82.9679484662575,
  17.4875082137668, 20.5702167389426, 82.712024280657,
  5.40970554857201, 8.79134279185671, 88.9936831196938,
  6.09295064194558, 8.06387216281591, 89.056632514162,
  5.61709971426515, 9.50248185025346, 89.6654486291233,
  25.7535267830301, 19.2334359260128, 64.770216108226,
  26.0079565087909, 19.7412325387341, 65.5932641716817,
  25.6590281577471, 19.8678366503821, 64.0030096622551,
  16.5245179406604, 22.8943615226475, 58.7480652039431,
  17.3731981484055, 23.4190831021884, 58.8144667773105,
  16.0006133499497, 22.9994762276609, 59.593331362394,
  29.8722390590099, 4.54557185855051, 77.0057774366252,
  29.7630235600963, 5.17029972264868, 76.2326105266915,
  30.8262045912729, 4.54990093094112, 77.3056624519002,
  18.8487549535899, 9.70456555572413, 90.7509036286674,
  18.5469642075298, 8.80013245831507, 91.0524382334867,
  19.7762992464489, 9.87458436429302, 91.0837026513786,
  19.366711239245, 17.2065828250213, 90.2749534484752,
  19.039610836322, 17.422399817874, 91.1949688570438,
  20.0833662828142, 17.8539783486618, 90.0155607259539,
  26.5880187412687, 27.31343560823, 87.0522454386332,
  26.9513037314795, 28.2213202891058, 86.8430340094077,
  26.9219522789022, 26.6568108176773, 86.3759819715767,
  26.2742170303863, 5.66116936215902, 64.0532788512959,
  25.9561757506851, 5.27035924415184, 64.9170596082413,
  26.5224162230315, 4.9237416337626, 63.4251088853135,
  20.9856609157503, 7.21554495516807, 80.5392195261055,
  21.3517806555451, 7.17059355951625, 79.6097381071618,
  20.486938115944, 8.07386422318441, 80.6598992804361,
  12.8543440016899, 22.2534467051544, 70.1769600383611,
  13.6649866059093, 21.9426127487843, 70.6731866194625,
  12.1844106682712, 21.5121953597377, 70.1352974449169,
  2.73033420884289, 14.8363519641376, 64.558446150329,
  2.20602218738525, 15.5340800104308, 64.0703145312232,
  2.76959813087039, 14.0026974002677, 64.0075574024261,
  5.15703240523968, 23.001054534012, 63.7578741664473,
  6.04415422721156, 22.5848353350978, 63.9573145120058,
  4.46881981486887, 22.2835617852101, 63.6503214543857,
  9.77441778449214, 24.9249146634177, 86.3288368611622,
  8.81062129624517, 24.9753282088711, 86.5906665838401,
  9.89939891076152, 24.1955862182959, 85.6561855865684,
  27.2889808803123, 17.0670124064079, 78.279454951147,
  28.1779348834514, 16.9820357763324, 78.7294991185839,
  27.2301977942992, 16.4072356818784, 77.5302959409443,
  24.2239843432531, 5.38518325249893, 61.6285468333364,
  23.7923897140394, 6.21120614347991, 61.2660385443148,
  23.6211748684286, 4.96408517106364, 62.3062614804212,
  30.3848583546072, 26.2586489514959, 71.9037202103254,
  30.8476015935219, 27.045712997834, 71.4958000198461,
  31.0604487943303, 25.6633544323666, 72.3386937649807,
  22.4398495865336, 9.08455069154483, 66.9855866188986,
  22.2370604739918, 9.30179525166694, 66.0307665432132,
  21.791946417454, 9.5602171087275, 67.5805344679251,
  12.0617892368447, 7.26749726591211, 71.7540320073584,
  12.2387803227197, 8.19905148061807, 71.4364144691394,
  11.2147642618007, 7.25174705526726, 72.2853517063311,
  8.54907483102683, 8.55347361000971, 77.695042041499,
  8.57008973241916, 9.36322195379451, 77.1086411601412,
  9.48450147198533, 8.25715647273027, 77.8878454479513,
  1.6235931447043, 27.8952838460825, 67.0749352409922,
  0.636297188042997, 27.8259859842555, 66.9319509750519,
  1.86622856197281, 28.8455140053836, 67.2703596474555,
  15.8163113983053, 19.6783238450262, 58.9687725371279,
  16.4632423391159, 19.7974403426503, 58.2155848992741,
  15.132839212949, 20.4077194028293, 58.9396539502576,
  3.27263287474541, 13.8808461229151, 57.7234787700489,
  3.46879991610443, 14.2310437512192, 56.8075747832606,
  3.74907088896175, 14.4389262686205, 58.4028559624678,
  16.8549054690612, 23.5349968197636, 84.1054354605056,
  16.6572861965815, 24.5036584163816, 84.2559058375969,
  17.7155707257689, 23.2965682494293, 84.5553322628332,
  19.6197140314437, 25.6110796041708, 63.8653528973999,
  19.3250785455813, 26.56129099976, 63.9667838303695,
  19.1898228557791, 25.2135023570288, 63.0547198672064,
  4.61863914718918, 26.7720053005414, 81.9295515165855,
  4.96265275552524, 27.6560120670878, 82.246074302463,
  5.36438697927219, 26.1057837082952, 81.9265580289095,
  16.5730737421074, 21.1954110530832, 79.6582035487382,
  15.8217828139471, 21.8204660728981, 79.4463824839965,
  16.6257263464945, 21.0607142862583, 80.6476905290761,
  25.836044088032, 22.8737714323097, 60.4645283344635,
  24.8872611448912, 22.6297352071175, 60.6651704227679,
  26.3379738317591, 22.0562189121239, 60.1822617776421,
  28.9099066077889, 16.6334846081712, 74.5798674591114,
  29.053656848548, 17.413704387349, 75.1886309307992,
  29.087638081652, 16.9103120780646, 73.6355274381916,
  9.73613103174843, 0.602955624704098, 74.9859563294286,
  9.90097090111286, -0.325231582149923, 75.3195673701639,
  9.38124479665329, 1.1670377421603, 75.731521299707,
  21.9365328346163, 9.53985372048664, 75.2623637942573,
  22.9013197407193, 9.72580331726969, 75.0763289231487,
  21.387398899227, 10.3330828350273, 74.9992298115621,
  4.29620838391507, 26.5779283212087, 77.4025857692409,
  4.74384912740246, 27.2608248070471, 77.9798813212762,
  3.55404507806965, 27.0096563125532, 76.8899410882519,
  23.5176012334238, 14.0772873239553, 73.8645332450093,
  23.4764565719361, 13.0824480993139, 73.9572803956172,
  23.3667332870952, 14.3294892115326, 72.9086916939806,
  7.16181035360007, 7.30557989109195, 70.2558093735299,
  6.81551823971639, 6.41053710144369, 70.5368434934525,
  7.97295284566903, 7.18452349954043, 69.683626528956,
  24.219061285879, 17.727608884064, 86.5620451182928,
  25.2141621773778, 17.7260664196274, 86.6608977183685,
  23.9135236723418, 18.6369945202181, 86.279796059002,
  2.87896785528346, 16.3712417636957, 81.1251478443668,
  2.49984657508605, 15.5485353051064, 81.5487291681962,
  3.86170666818207, 16.4159766175387, 81.3046561129069,
  25.8244282846279, 4.71691754966296, 66.9394768991763,
  25.650093480646, 4.36798509328993, 67.860266515218,
  26.5598127715458, 5.39372972279423, 66.9731657504748,
  19.1674180668794, 7.14654155217814, 73.1818818111505,
  20.1334679868321, 6.97060113653701, 72.9926926933256,
  19.0869603167298, 7.90882066656463, 73.8241100433321,
  30.6879805314817, 29.9534725088829, 74.8811160482269,
  30.5042813147455, 30.7003430993689, 75.5202083098274,
  30.4772015180663, 29.0799108431534, 75.3198212153625,
  18.4756618005605, 8.17128439642982, 77.9344451012673,
  18.9575422426228, 7.47744917439911, 77.3992965945633,
  19.0086880324303, 9.01736249825375, 77.9403511788706,
  18.6069963618542, 28.0915383817735, 63.1146979245993,
  17.8148429860048, 27.4832131630584, 63.0653678383878,
  18.3017061558382, 29.0198428389639, 63.3269447735067,
  1.94290819467519, 24.3802856748939, 60.9979171954008,
  1.50126282850073, 24.4483474456401, 61.8925215581778,
  2.16063660443185, 25.2970473230953, 60.6630404718564,
  11.9636453331041, 28.1935207013298, 71.9335608957181,
  11.8925798906395, 28.8992921692804, 71.2286947113156,
  12.5013886775999, 28.5420621162808, 72.7012528766027,
  16.6128124883941, 1.25504645916675, 67.0859718872798,
  17.5415568009892, 1.37623235783099, 66.7356178095426,
  16.0468995659781, 2.03030926427532, 66.8054185995468,
  30.3601847887309, 13.0926247166845, 81.1428824100985,
  30.5739973201611, 12.5775604533514, 80.3128263842541,
  29.3942778433686, 13.3513971054328, 81.135096286398,
  24.2423677061974, 16.838798610776, 62.9129942952598,
  24.0535434037672, 15.8783098597411, 62.7085273249512,
  24.3038202476895, 16.9629490863009, 63.9033529396767,
  4.90841520662218, 4.65095313811927, 76.6220385260798,
  4.69163572021761, 3.72027530019046, 76.3273430624868,
  5.75589435475888, 4.95049375852862, 76.1837982835207,
  24.1007555407931, 11.4482719483529, 77.7479956312134,
  23.7842294977426, 12.2559391462556, 78.2454742352789,
  25.0687027520565, 11.2931995646584, 77.9455576519124,
  23.7745359204124, 14.8629602170892, 55.2480395861575,
  22.9714832070849, 14.5542101223143, 54.7383536842592,
  24.6039415715059, 14.5898283868581, 54.7607149825834,
  21.9647490996366, 6.89344562278065, 71.5045495030607,
  21.9381204700959, 7.23002202039595, 72.4458290814311,
  22.767452077093, 7.26690357536815, 71.0395795173286,
  4.92732158300977, 3.53583160302578, 67.8782972552745,
  5.03249222555121, 4.44525615890999, 68.2806479892148,
  4.63970449798518, 2.88975248967665, 68.5853037557368,
  2.1170565540641, 30.1458137952421, 77.1815640825334,
  1.77277063168497, 30.8646375488939, 76.5776107607962,
  1.98131973759965, 29.254172064686, 76.7496491129074,
  27.2962528000376, 18.043176680852, 70.1705944919438,
  26.8480254972065, 18.3671488776126, 69.3374472656249,
  26.6551487539588, 18.0961773093569, 70.936216157964,
  6.42482237222944, 9.42218986859551, 57.7235578315522,
  7.02002613714363, 10.1935021489327, 57.9489682226904,
  6.97014362275934, 8.58591684356178, 57.6663550228672,
  22.395224746184, 15.9392920283841, 88.1007684861938,
  23.3552671025115, 16.1894539169169, 87.9753184818779,
  21.8248457219816, 16.7570469401601, 88.0236667805303,
  6.27493157956827, 20.4968224392683, 87.4839004625112,
  5.94206717123192, 19.5699071764934, 87.3106105860099,
  6.75030368438692, 20.8373944202383, 86.6727086924972,
  20.7062850608531, 22.2662409632249, 90.5103194326296,
  21.5691175677128, 22.6501167551985, 90.8391954600972,
  20.8493784632813, 21.3174061776859, 90.2288290634646,
  1.66533919704551, 19.5667689778007, 56.7311116735154,
  2.47288389139342, 19.7076249511766, 57.3038517204781,
  1.87857240352453, 19.8173990041816, 55.786804419741,
  24.0540716308857, 6.81350583687449, 81.5741930696864,
  24.1738998651763, 7.80447565602177, 81.5140265357493,
  23.079119086212, 6.5931727364811, 81.5438473862155,
  18.2215857684036, 6.07250723792459, 84.0487324702578,
  17.8541060782392, 5.61899804340905, 83.2367668996783,
  18.5643961099985, 6.97794532156613, 83.7984067896192,
  24.1317413990209, 13.31810478971, 79.6544460105787,
  23.3466078536541, 13.4441822583006, 80.2608038157182,
  24.7818159454388, 14.0656023785099, 79.791012620106,
  5.93809759005122, 11.9526689216871, 89.1393944945318,
  4.9759103175326, 12.1184701441836, 88.9232796935074,
  6.36209546684536, 12.8043170584681, 89.4474874214085,
  21.7400649017519, 11.9161517619281, 84.6962590114602,
  21.6749001036854, 11.7475034123791, 83.7127391675895,
  21.7038645737563, 11.0455292719807, 85.1868770056785,
  18.8444104670216, 22.9088219576882, 80.5840176392178,
  19.4617186861967, 22.9092358304467, 79.7972963472419,
  18.2003791325671, 22.1482337428623, 80.5019858910422,
  30.8903882110329, 0.145051993747046, 80.6716564387381,
  30.9038672140443, 1.14453517312175, 80.7008401777868,
  30.0386334326968, -0.188769437657299, 81.0754844337022,
  27.8898815506893, 2.05395958199036, 81.7873802613549,
  26.9506501853886, 2.39649848947443, 81.7647630268877,
  28.2610057743026, 2.03711035540996, 80.8589499116727,
  30.116432245975, 1.60370199310817, 76.2499059420257,
  29.2219139038979, 1.18419321805494, 76.404338203361,
  30.0834763091856, 2.56685012730636, 76.5168508386258,
  8.03066568251899, 1.89319642576839, 70.5116842616842,
  7.85675394417499, 1.57249577739671, 71.4427620250316,
  7.97814104036874, 1.12138206538665, 69.8780094593797,
  26.2633301919967, 10.0085867878419, 82.339731106636,
  26.1411695730238, 9.04610696426417, 82.5820312766275,
  27.2376879927044, 10.2334260509038, 82.3483440031134,
  10.4890313277414, 1.43888890974364, 89.1148612060008,
  11.1150016100462, 2.21499231531156, 89.1911809907036,
  10.5687241210899, 1.03470666227709, 88.2036610251837,
  13.3516269857767, 2.28716033969797, 91.5193847232491,
  12.5106836814763, 1.7463462146064, 91.5010969936512,
  13.1743621595639, 3.16406715520137, 91.9661638838099,
  0.166368074561163, 9.7566207119224, 87.0726087745983,
  0.601958927522787, 9.19598215804622, 87.7768424153197,
  0.866893076224365, 10.2596889512456, 86.5664595193098,
  22.9548807939073, 20.5008237283526, 69.2237203479619,
  23.8032319210728, 20.9966068079695, 69.0379799296287,
  23.0490131540955, 19.9868101002094, 70.0763217136942,
  7.02476593377206, 6.16483684553301, 88.7488323490492,
  7.43044232836382, 5.59027448145209, 89.4596802601053,
  6.80584725759604, 5.60324350599949, 87.9509053259369,
  7.81700033592767, 30.6858802598114, 69.138066424975,
  8.54191533934292, 30.2849589345216, 68.577923292596,
  7.19350990289592, 29.9654971681101, 69.4418885458101,
  2.53007490296129, 2.45038749246476, 78.8984560762361,
  3.47747639219886, 2.76111186767352, 78.9751423256004,
  2.51333442108143, 1.5172888811107, 78.5392253178711,
  11.3725715003207, 0.472555904897302, 86.0008414771305,
  10.5166216561026, 0.0115614309251929, 85.7666749569999,
  12.1302879711763, -0.176419070788703, 85.9323051310979,
  16.6861844946712, 22.631672942929, 74.2485391025022,
  15.8592533579692, 22.2797365839298, 74.6870886371811,
  17.4176031116026, 21.9538970247599, 74.3236830414202,
  27.7634979833891, 14.570717172864, 63.2628089474552,
  27.2431982996886, 14.9050012473505, 62.4769702892779,
  28.3346578097704, 15.3084702420557, 63.6226656712026,
  15.183416070144, 0.851285613086289, 63.3080578139254,
  14.8844582946418, 1.79978577131015, 63.4128036888613,
  14.6817527557158, 0.270884319187148, 63.9495157291445,
  10.9507047495709, 21.1303032800393, 62.3326197598132,
  11.5848816649117, 21.3258813949643, 61.5845764181469,
  11.3154541064509, 20.3867604729658, 62.8930677954997,
  27.1097408998614, 15.58757878719, 66.6608447760369,
  27.0341899739698, 14.597328091581, 66.5438164997843,
  27.6530753055823, 15.9710131585698, 65.914007573961,
  2.9450022561875, 30.2910698711224, 70.4275883641429,
  3.38346620055625, 31.1324353197196, 70.7435844897448,
  3.43511596141832, 29.5010941712636, 70.7959997504729,
  6.01031130886418, 3.79403296453967, 86.7741835816949,
  6.65100134973178, 4.13336860289031, 86.0854400909248,
  6.49270372314546, 3.19162485655395, 87.4101097016782,
  22.0904373580422, 23.8359256227768, 73.6057288837496,
  21.8844018471069, 23.8621223031421, 72.6275350879343,
  22.5465527343353, 22.9740427477774, 73.8273517013741,
  13.8607755965073, 20.0894079273231, 78.9872903674932,
  14.1120137300996, 21.0442965705077, 79.1456162319185,
  12.8653045693308, 19.997937415812, 79.0131859187737,
  16.2154218635527, 25.5004224847832, 67.3282333341707,
  15.4330844242, 25.3311310323645, 66.728826514786,
  17.0614744225441, 25.2828672976391, 66.8415457465224,
  29.1831581053827, 2.76422214605429, 87.7626658665952,
  28.2534926669064, 3.11406204938825, 87.8781397360983,
  29.146456824335, 1.83623940376439, 87.3918545318418,
  24.9159762227763, 0.770660763755038, 64.1553435680596,
  25.6906255939528, 0.916792132901148, 64.7706190955165,
  24.9679428605048, -0.149224022969518, 63.7666130087825,
  14.0669075723676, 0.128732211813464, 70.6613552501344,
  13.7280295299191, 1.03302446774159, 70.4017070492651,
  13.8607110523542, -0.0404355796530567, 71.6251318079862,
  28.8680527402424, 26.7270088842812, 89.0738295763413,
  27.9946368440169, 27.1522884882663, 88.8365914456481,
  28.8621400142911, 25.7697427943144, 88.7846813917171,
  15.0766567998791, 22.7467862105509, 65.5263941509143,
  16.0755872080672, 22.7304947997841, 65.4831202611834,
  14.7698344096963, 22.2456375777119, 66.3355357137363,
  14.9349755242545, 29.7072955301061, 80.3002794413756,
  15.0976818129665, 30.6527442487668, 80.5825087523914,
  13.9882812531508, 29.4570758203696, 80.5031588487061,
  24.4038328766031, 18.4293830067953, 83.1170376492031,
  25.3280003842809, 18.5250409024292, 83.4868537991419,
  23.9812712989421, 17.6014562333385, 83.485790914786,
  4.19162478831251, 15.934550183155, 76.0630505366538,
  4.03113555161289, 15.6433949816396, 77.0061686912527,
  3.4094225965113, 16.4679882155131, 75.7411754105951,
  5.6705087696452, 28.9828650045771, 66.9217409010871,
  6.18915671015347, 29.8059307015663, 66.6902950710398,
  5.23189933447548, 28.622719732001, 66.0983836602607,
  24.1664792299012, 17.9956729528508, 68.3845822941289,
  24.3203560165255, 17.9168771025739, 67.3996390731678,
  23.5856263115196, 18.788551772269, 68.5688458687322,
  15.8936053948099, 3.95846819086621, 72.0273488063786,
  16.7024922860343, 3.59122435201527, 72.4865153992741,
  15.4004115261203, 3.21503933616159, 71.5756040267966,
  27.3440813247829, 24.1903922359058, 83.0543497294734,
  28.2950646007469, 24.179933213379, 82.745284335609,
  26.736415485745, 24.0898965212789, 82.2665408443952,
  24.7611201491648, 29.5738131396358, 62.202811871017,
  24.9460420271193, 28.6318064732249, 61.9227630547524,
  23.8231778499296, 29.8170429140787, 61.9556206087728,
  1.64452954088434, 1.00217715587739, 62.2816297809042,
  2.59730480149716, 1.02662764298987, 61.9789393838908,
  1.47812400584428, 0.157813932704087, 62.7909037202143,
  12.6772453189116, 6.97804454073839, 86.1783490334373,
  13.1330116999446, 6.1195875975464, 86.4135695312805,
  13.3175106648202, 7.57321248424655, 85.6927201567744,
  15.4171953939985, 30.5530311402007, 83.9926202398795,
  15.1541341903573, 30.2110349255893, 83.0904908742504,
  16.095408910583, 31.2804940544917, 83.8885811402425,
  3.40019002143191, 9.56557456683268, 56.9951206071186,
  4.18318491472822, 10.1844309223752, 56.9323845865521,
  2.56746053461956, 10.09646095399, 57.1523505206982,
  11.60119633304, 15.567263911613, 71.459457120607,
  10.6093927086531, 15.6080059763788, 71.5805589571397,
  11.8221426788832, 15.6520166695222, 70.487860659989,
  25.138739244138, 2.74142745943194, 81.4794859598387,
  25.1057017104965, 3.5825910802618, 80.9397153749017,
  24.3416714241982, 2.17664606147152, 81.2656990029533,
  28.6109309338096, 13.620942957355, 78.0220150595283,
  29.1575603735515, 14.3816065894852, 78.3721394579383,
  28.0398519855848, 13.9410421926367, 77.2661014967008,
  7.79100308767522, 9.85896009627108, 65.2564981823977,
  7.03346060380308, 9.4907095712181, 65.7954981229609,
  7.82406873750662, 10.8526756474632, 65.363437726628,
  25.9245250473773, 25.5415374068229, 68.5521522788093,
  26.0332030138325, 25.2576451212648, 69.5048297005045,
  25.6191601566969, 26.493252916035, 68.5206900305601,
  6.72431432195721, 25.3002039953381, 65.2538369992484,
  6.14387713732517, 24.5212891712608, 65.0163830636546,
  7.29226447860729, 25.544536928456, 64.4678764166775,
  14.7649765012297, 6.13728295455788, 73.0207188438986,
  13.9305406971151, 6.51537586901677, 72.6197666811067,
  15.1731203303191, 5.48216020109078, 72.3849258015759,
  21.2888055674566, 7.19069577914694, 87.0113464266125,
  20.3237054160958, 6.93028789589487, 86.9836077859904,
  21.847537307407, 6.43690063471106, 86.6654971487517,
  24.0905343761394, 21.8030799780815, 74.0879194880122,
  24.8115154043346, 21.9001595286969, 74.7740404087214,
  23.5194040642973, 21.0139349431091, 74.313884708065,
  20.4520122754998, 21.7661479685705, 82.8699479553691,
  21.2544313163053, 21.3786977135406, 82.4160691358259,
  20.0899636510181, 22.5196135839706, 82.3211216076773,
  0.738046350484638, 30.5434072894315, 84.3224906818956,
  1.46160292211647, 30.4968990844383, 85.0111871858193,
  0.788614363673695, 29.738684793347, 83.7309971651622,
  3.12630738020732, 6.77963136016002, 56.5702189099977,
  2.25904543209921, 6.74252887780153, 56.0737512683869,
  3.39081137380424, 7.73408389887742, 56.7082695844154,
  0.469297354323308, 18.0365469317123, 58.6713035820493,
  0.700796692800825, 18.4798253305136, 57.8053288032938,
  0.718788270153192, 17.0691501504684, 58.6277404031323,
  17.1925658378026, 0.878358514334352, 72.1907376435286,
  17.9439705181828, 0.473030774289235, 72.7114106978081,
  16.4327681632908, 1.08437667629009, 72.80739314764,
  3.20025135568273, 7.75453992925218, 71.3805275113987,
  3.80134813402226, 8.54533135914173, 71.4959899619316,
  3.18993380163085, 7.21767594797523, 72.2241332330992,
  0.735213906732909, 17.128046453597, 86.5350124174195,
  1.25719720542424, 16.370311179923, 86.1433867148443,
  1.30773025639821, 17.9474307918219, 86.5638972860826,
  12.3610913570175, 25.2462073795762, 78.6357383834083,
  12.9042324697418, 25.79212054597, 77.9977912489008,
  12.6746344274709, 24.2969089230455, 78.6128651807633,
  15.6886582275229, 13.0711790470704, 89.0027178844031,
  14.8328741678985, 12.5879399134603, 89.1874165120114,
  16.3858578468307, 12.7759879747012, 89.6559980093347,
  12.4944040574907, 19.0152940445714, 63.3514084149489,
  12.1563653095776, 18.599531313554, 64.1957253912121,
  12.6043332631623, 18.308509572416, 62.6525727549683,
  11.1135837469522, 24.0554851270251, 68.7762030885072,
  11.4334225412399, 24.9715309991479, 69.0182012410524,
  11.7266448881836, 23.3725925759992, 69.1734609403685,
  -0.0772392704062469, 27.4353025179799, 82.4049337845804,
  0.766358775771906, 27.7312652974884, 82.8529833015202,
  -0.10460215972362, 27.797477429948, 81.4732253508796,
  14.9781539730548, 8.74088085635784, 74.9823153326151,
  15.3496300221973, 7.83966710727429, 74.7591129057103,
  15.6741562428459, 9.28026728337931, 75.4562806507457,
  18.880459285278, 8.94118793349081, 83.4055419928801,
  18.6772859891657, 9.03595759979248, 82.4309962925171,
  19.4661782525706, 9.69672885531625, 83.6989550239486,
  17.4132391034567, 17.6277773445568, 75.4867013738254,
  17.7026722850756, 18.3913484241772, 74.9094772927744,
  16.8967287767104, 17.977769687719, 76.2681887007171,
  25.8302321059148, 18.7588580525134, 74.9421962732359,
  26.7342870882716, 19.1753553064564, 75.0381891184583,
  25.2608955601669, 19.0142121668735, 75.7236373611979,
  9.11766682443479, 8.15517812870724, 88.6681313130586,
  9.49816900628325, 8.43927720619635, 87.7880711993286,
  8.3941345019346, 7.48170868064621, 88.5166721409169,
  10.2446892427203, 22.5751996882099, 84.7540114382166,
  10.5220641268151, 21.8505891297732, 85.3848859996593,
  10.9225498382447, 22.6587751767197, 84.0235868009297,
  19.0247065260408, 16.102902212079, 77.5138349851077,
  18.7432130647897, 16.8402042484394, 76.8997119205257,
  18.2981067955253, 15.4179257383847, 77.5673145335359,
  18.3551643898299, 27.4773603213472, 68.8428028799203,
  18.597525584122, 26.626517579865, 69.3089870503598,
  17.4154148026274, 27.7285261717695, 69.074721893661,
  13.6146153714833, 10.2337768848244, 79.7501645763146,
  12.8573390753915, 9.8580702804942, 79.2159575388841,
  14.4173811818582, 9.64603314282889, 79.6495447599849,
  21.9826064413617, 24.4144685217718, 70.7626615745277,
  21.3288458580747, 24.2271260487041, 70.0295177294843,
  22.5132061305197, 25.2310896303073, 70.5355185910136,
  21.4075719467239, 19.6363357070858, 89.8335232400556,
  22.237986231081, 19.2248557835157, 90.2091512326685,
  21.4526536676352, 19.6255376929688, 88.8345982972642,
  10.8122473134119, 6.33555115674085, 75.8493801010743,
  10.9110448839613, 5.38910220283399, 75.5420148172472,
  10.455179149114, 6.89371559428385, 75.1004109517049,
  10.9359854614916, 3.77176487181715, 72.162116821587,
  10.2245010123664, 3.74977814038729, 72.864474609537,
  11.4511484262534, 4.62565837445907, 72.2360965883056,
  26.3766009309779, 24.7692512925637, 64.2805064845166,
  26.5442592457577, 25.6846668708923, 63.9145761517502,
  25.4692165595686, 24.7388659332803, 64.699708503194,
  11.6290703874072, 3.20914735475428, 59.0317750190396,
  11.6929462875327, 2.27171523101082, 59.374033521866,
  12.5203531645618, 3.65521656271161, 59.1132444787159,
  23.1873308928478, 4.80981575199793, 86.2585706474669,
  23.8508002489546, 5.20862132187066, 86.8916287261183,
  23.6712220841178, 4.36893336859123, 85.5026129508907,
  20.1641425110273, 16.2690290299947, 59.1044205798975,
  20.4775486899892, 16.7500102566702, 58.2856204659659,
  19.4685567215211, 16.8180615578714, 59.5678034591349,
  0.303248932639976, 25.5407724195513, 79.4890378531551,
  0.192357730674553, 26.5224718014946, 79.6438586037634,
  1.17153586832395, 25.2373971606529, 79.8815187439114,
  2.73663756786986, 7.90228738109625, 83.1716394374222,
  2.95870119488575, 7.65440467986931, 82.2286431956539,
  3.5134356130769, 7.68892951058447, 83.7641453159189,
  10.705598792232, 9.34647665629995, 64.9981169138271,
  9.7434182066261, 9.50099810283989, 64.7737697648762,
  11.2207692014865, 9.1772084486672, 64.1579099611581,
  4.56713836967944, 0.348358609756652, 82.0469830531167,
  3.83693494450867, 0.808212185139585, 82.5522925098622,
  5.28705611237936, 0.0686402480260995, 82.6821807245991,
  15.7133492898058, 24.6116990792286, 81.0474353334529,
  16.5446493791526, 24.6117045973496, 81.6032591917223,
  15.092601551276, 25.3234942062066, 81.3760992078301,
  22.7464243116745, 12.8094287408779, 62.5936287342701,
  22.1518035151735, 13.5830593519795, 62.3747182824065,
  22.3206753647323, 11.9617494081051, 62.2771203094732,
  3.77774840362722, 27.4659030172618, 65.2816943927056,
  3.87381591264273, 26.4749951188424, 65.1875000693016,
  2.93427103035222, 27.6734345061593, 65.7771503462365,
  14.1446116290201, 17.3127113730172, 69.4720318809696,
  13.7619217050536, 18.2365815041555, 69.4685101079787,
  14.2176522019945, 16.9857451126543, 70.4142410611859,
  9.3428160215384, 28.0584336181638, 64.2628763272423,
  9.83922660414996, 27.4940388665106, 64.9224482321758,
  9.97301510252662, 28.7101649381253, 63.8408628145406,
  2.52190878537472, 3.33642340434688, 63.8126498298161,
  2.23626063087793, 4.29414399126654, 63.7783510073461,
  1.89231707781308, 2.7811223126377, 63.2692761284685,
  16.7731249517977, 11.728460712262, 79.9821859379061,
  16.7668188486675, 12.4172843252473, 80.7070874920894,
  16.0860345163153, 11.9622130364988, 79.2942422015566,
  0.563858623903612, 7.33266697514936, 85.0212983649078,
  1.25867768975367, 7.78030259767424, 84.4584051111038,
  0.00435061039287831, 8.0265215506002, 85.4746377641918,
  27.3195159455287, 19.9291785289545, 83.4743823070815,
  27.9874929178548, 19.2157645645325, 83.686154070567,
  27.4637375495515, 20.7113833279729, 84.0804811285006,
  17.1943068799329, 4.81714571239833, 64.2119892732277,
  17.5507175707458, 5.01788949503843, 65.1244986447991,
  17.4942793627608, 3.90582835212952, 63.9300013684893,
  13.856467864978, 25.3581396713841, 65.8500668249604,
  14.2602525178321, 24.4433055665374, 65.8440240831361,
  13.1101425807603, 25.3974962093171, 65.1856500633871,
  5.7724916672564, 25.6290507644077, 92.2414108027986,
  6.31831604388916, 26.0966153027475, 92.9367230724736,
  5.59572469417205, 24.6889586080992, 92.5329243957473,
  24.5624048461017, 1.79260903470404, 61.0573538196771,
  24.4719611089922, 1.15655944289362, 61.8236832835342,
  24.0006524878374, 1.4757961546159, 60.2931130938618,
  19.9563086862223, 20.249140350627, 62.6949363551881,
  20.4708518203667, 20.0787301319886, 61.854575884623,
  20.5886062908957, 20.3033323612099, 63.4677642565434,
  12.1400224159606, 19.3335924651582, 69.5300070299435,
  11.4524675169122, 19.1468253193601, 70.2317094555093,
  11.8099997822187, 19.0064812082328, 68.644522254913,
  29.0221925893855, 6.88521620074409, 75.2140292186945,
  28.3411522737581, 6.32053499724141, 74.747854115433,
  28.6105095545041, 7.75937074714311, 75.4716547372302,
  14.419628660123, 21.3779872884224, 63.1925280906438,
  14.5612340230354, 21.9175292025458, 64.0224934176897,
  13.7855613093729, 20.6292540924441, 63.3858081877905,
  17.3426068552552, 11.1255045088666, 60.9164272705842,
  17.3658089609979, 11.0044798298599, 59.9240489710631,
  17.9239108591774, 11.898111329737, 61.1717003701629,
  30.0534875877028, 22.8124167220277, 62.7176433830929,
  29.2211000243716, 23.1930296300335, 62.3148223823111,
  30.5544470294004, 23.5355126549115, 63.1932187289856,
  0.78679514085643, 29.3188668594949, 91.9406277421809,
  0.267129105770296, 30.065126732125, 92.3566126150789,
  0.886472760285149, 29.4881552879394, 90.960114713109,
  21.7541196439666, 11.3741029146828, 81.935528321062,
  21.0457155300906, 10.902849251309, 81.4100917442991,
  21.8016009109524, 12.3306919037473, 81.6479817417292,
  14.4450208643252, 12.3400625524907, 71.135671264773,
  15.0505702016849, 13.1329760038832, 71.0678608037503,
  14.3176586757629, 11.9393317330844, 70.2283710480297,
  12.7828282517906, 15.7165574505468, 79.802343399969,
  11.8858271729837, 15.2897433260014, 79.9173162998533,
  13.2597556013025, 15.7319721329868, 80.681150939111,
  16.3096936979351, 14.5839631883326, 77.6811806905433,
  15.8362844230205, 13.7142009487975, 77.8204548988649,
  15.6477553036107, 15.3327953951736, 77.7141638395278,
  5.21658456505446, 18.7993034320448, 61.7192844963325,
  4.94339749148739, 18.3696085825093, 60.8586270969461,
  6.21365846386388, 18.7893536571453, 61.7950779148623,
  17.6905398642856, 2.14434628396043, 69.6221254582471,
  17.4266020100482, 1.72133222818474, 70.488956420844,
  17.3051034242531, 1.61874630357367, 68.8637169856464,
  9.02214555828264, 16.379161481469, 64.9482710122352,
  8.27616352979973, 16.1494847426538, 65.5733785300493,
  8.88475024176084, 15.9069614438564, 64.0775531179224,
  11.7719968088095, 12.8278112636116, 84.2702823577757,
  12.1972655730795, 12.5857492621667, 83.398185765882,
  11.5483413406059, 13.8024759581725, 84.2729214332326,
  15.4699736360891, 7.206848999803, 61.2304070970787,
  16.1274659117187, 7.53171668432857, 60.5505799903534,
  15.949634132557, 6.68294372507092, 61.9342885297334,
  15.0367404170067, 2.19822093255067, 74.4844927198854,
  14.1854838136842, 2.28726687286337, 73.9673534583575,
  15.3202352213903, 3.09759604182139, 74.8172916211934,
  26.8569676481474, 20.4973255303882, 80.7045796515497,
  27.747934373736, 20.9469783156755, 80.6414079286251,
  26.7552400154825, 20.0847305557024, 81.6097961315237,
  26.1008981003931, 10.51815445277, 65.4606452624569,
  27.0579225701749, 10.4535488306875, 65.1779258293888,
  25.6391060195541, 11.2185853044559, 64.9164534800115,
  5.06154696180431, 14.8440718047214, 68.4649541366473,
  4.79099450596751, 13.881588677062, 68.4856325701399,
  4.32808298624566, 15.3878222845426, 68.0570742373487,
  3.13141467573311, 9.36269303487744, 59.9182813492521,
  3.27853793330906, 9.60246662960636, 58.9586650872229,
  3.9937258455523, 9.056016350032, 60.3212315414313,
  9.31638432096348, 26.174473232586, 66.3345608910992,
  9.8379359672276, 25.3599262445126, 66.5885236531328,
  8.38652855704769, 25.9089284400765, 66.0798959710893,
  16.6845690838585, 26.2900930691797, 62.4608134029078,
  17.4020284701319, 25.5994179598561, 62.3701496151581,
  16.4630856374358, 26.6610413075537, 61.5589583771925,
  16.2004795915264, 18.8485515393659, 77.5338230518666,
  17.1287586056991, 19.1399477120421, 77.7648778990264,
  15.5630168042697, 19.1861484664236, 78.2264048229985,
  29.1128643138476, 13.0148599122832, 61.3846624675076,
  28.6679723885269, 13.5496425255515, 62.1030486667976,
  28.4842247527758, 12.3100051188541, 61.0560410707066,
  22.7756176814371, 20.078110008755, 81.3935234357187,
  23.3687091895868, 19.6221890845401, 82.057133693192,
  22.1428208129551, 19.4118346813224, 80.9990043470882,
  30.5294894084837, 9.3094098936348, 77.2160499858063,
  29.6823275494419, 9.18571447396296, 77.732786115506,
  31.0665369865772, 8.46652727330204, 77.2496474143535,
  28.7223804558085, 4.90859509434129, 68.3461709773937,
  28.2845580406428, 5.7925059603043, 68.1818143109303,
  28.7854084289493, 4.74577646492118, 69.3308118096344,
  11.3747991816099, 28.1195627487842, 76.3436302820508,
  11.3258996914394, 28.9001421009168, 76.9667712892757,
  12.1789248163813, 27.5672948665825, 76.5635897096552,
  6.74728973047572, 19.4295130254928, 79.2757683160926,
  6.8550700209981, 19.0922321909261, 80.2109822208272,
  5.84477139604725, 19.8480357198743, 79.1742823056869,
  11.293519704755, 17.5735834851141, 57.8122648058475,
  11.9898377951419, 18.2815444868239, 57.6942294846165,
  10.8646432446428, 17.3775311080048, 56.9304323685946,
  3.89515225402209, 11.0052570864147, 73.9368571851991,
  3.30463790205431, 10.3519103149568, 74.4105984609453,
  3.96325846100627, 11.8447743561037, 74.4759047698001,
  17.1566246832792, 30.4292915518916, 64.2383599500605,
  16.3442404011024, 30.9512264844838, 63.9783297514067,
  17.00725326688, 30.0024858527239, 65.1302820739709,
  8.64874710681167, 23.3177053239133, 81.6072472694255,
  8.7370421070927, 22.7164154633658, 80.813109689073,
  8.79228116070458, 22.7886032009455, 82.4435778971344,
  6.21633613868071, 4.12062824010044, 61.4544439565532,
  5.57323536023534, 4.82611533707282, 61.7522850967076,
  5.73979943439415, 3.24450021058066, 61.3815574327131,
  14.1750046302938, 15.4182092608363, 64.3065099956581,
  14.3093993063048, 15.6295473489824, 65.2746392657241,
  13.2268118266588, 15.1391071605171, 64.154745623251,
  27.6263852651903, 12.8972733127905, 89.4666928865219,
  28.3833951738519, 12.2591196787029, 89.3263506708883,
  27.9403277421083, 13.6710470166046, 90.016887739708,
  4.38070338497273, 24.1224915172136, 86.2422932492996,
  4.24902880278626, 24.894112794781, 86.8645973617809,
  3.92470925000375, 23.3135026090624, 86.613246474602,
  26.0684011517368, 2.80980316144841, 74.3559674777758,
  25.5844231101906, 2.35254747694834, 73.6098558947713,
  25.6074075904416, 2.61432551730148, 75.221573292846,
  28.7677080059602, 17.5641575066468, 57.838907121552,
  28.7369080920071, 17.5715885395346, 56.8394091750555,
  29.6398695540037, 17.9430678389653, 58.1483601780512,
  23.0796714951559, 25.6417877295918, 75.7173893063918,
  23.1904016223429, 25.0896527961556, 74.8910202277034,
  22.1974197012635, 25.4353455865667, 76.1404890744807,
  11.2303917819326, 20.4961176452481, 80.4556619652605,
  11.5568984797278, 21.1659910780912, 81.1224924986541,
  10.3380970536077, 20.7815738300516, 80.1059122199268,
  12.089717566403, 22.9237586495025, 82.8407463930558,
  12.4366715196158, 23.8499792685312, 82.6933071878355,
  12.8579855732163, 22.2960487625644, 82.9662237517601,
  23.6124126534911, 26.6172228607473, 63.0510363066158,
  24.2405393597326, 27.0127320544437, 62.3809398071415,
  24.0342636269851, 26.6400787849855, 63.9574133599934,
  22.1602344403733, 9.4361032157042, 64.2516435041622,
  23.1251604677759, 9.409203708298, 63.9905033537787,
  21.7142590285591, 8.58730052061424, 63.9676718209521,
  28.1296348570214, 15.6261725237146, 69.1967882250203,
  27.8367755433991, 16.3913988632166, 69.77007878988,
  27.9592728616068, 15.8451282705796, 68.2360410306798,
  9.57081296417908, 16.2949781585425, 87.9946267280392,
  10.5389684192643, 16.5188628279962, 87.8825969571193,
  9.47774589831772, 15.3287378726351, 88.2348729166489,
  3.63045681880746, 20.4114602336706, 79.4530873566024,
  3.7508200384651, 21.341872517037, 79.7992747022904,
  3.27503620232089, 19.8275806901534, 80.1829920517773,
  5.09286142107234, 11.5952149042319, 66.5084062104905,
  5.23710962895558, 12.2527042129384, 65.7688791565843,
  4.67345269803607, 10.7656251244914, 66.1397910719093,
  26.965579958154, 26.3640465017385, 75.555471796212,
  27.1167182317238, 25.4817912894781, 76.0013226263129,
  27.2949199682173, 26.3216190467216, 74.6122141066953,
  5.73102424652159, 8.89469274863307, 60.7859502226271,
  6.36494550127766, 8.64683453130873, 60.0533451810983,
  6.12266519063055, 8.63349841138399, 61.6682171261695,
  5.82627425541259, 15.015841660263, 71.5881279471903,
  6.53222211129373, 14.9553327027733, 70.8824535953535,
  5.2205302568128, 15.7860471915149, 71.3884841449088,
  22.5793069938178, 19.3564812584913, 74.7593459031843,
  22.6937174229173, 18.7349911214983, 73.9843231529804,
  22.9232191321979, 18.9196253473809, 75.5905386329425,
  2.29715155909143, 17.6010019920919, 68.9666603639119,
  1.42275558606883, 17.1577154085875, 69.1639639047997,
  2.71894663080374, 17.1667240035652, 68.1707385422734,
  4.6208078269837, 7.06751636205145, 84.9378355076017,
  4.73141387908902, 7.83481659079865, 85.5695131628992,
  4.27722552726491, 6.2718786905716, 85.4367462200966,
  25.6888839440747, 7.38441586743781, 76.3743051661495,
  26.1984644900447, 8.15482147202665, 75.9911565375639,
  25.223785765079, 7.67520468556776, 77.210442443841,
  20.4415592379443, 30.7422462884397, 66.3600073139487,
  20.1828905187504, 31.7033738285286, 66.456569964043,
  19.6340927031352, 30.2018818944632, 66.1233554242756,
  2.23363571344491, 19.6431846461886, 77.2923958721747,
  2.67088114469103, 19.8111521986536, 76.4088782808539,
  2.89952372690148, 19.781467652241, 78.0255199842948,
  5.2260121334013, 29.9352039177942, 88.9518108584574,
  5.76985452753253, 29.6452008700759, 89.739296529857,
  5.83427575002738, 30.2656259023374, 88.2301206999963,
  17.0631706534525, 14.2927056173404, 86.7894731882051,
  16.7699474371078, 14.0475974760724, 87.7135630888535,
  16.4575003010609, 13.8598964647733, 86.1217609285543,
  11.5835800532373, 8.86580739942242, 62.3249813879837,
  11.5143088473417, 7.86994973534487, 62.3838797150549,
  12.5066778630752, 9.11922050300863, 62.0357198585623,
  5.31663363052077, 22.7751961206662, 83.9260339537635,
  4.9999234637745, 23.1200942731116, 84.809628846641,
  6.13900893168689, 22.2221100241735, 84.0594304825732,
  21.7777855537575, 24.684454915959, 65.7912833344431,
  21.2499551184248, 23.8363132308028, 65.8365681380412,
  21.6862338122722, 25.0858011489407, 64.8799439465625,
  18.6225424992281, 3.924631355549, 92.4675335260541,
  17.6555198217852, 3.67504221006634, 92.518252356565,
  18.70477347834, 4.90214566113395, 92.2733587376518,
  6.04717395642258, 20.9195487788, 74.6726912841008,
  6.4022854451451, 21.4564903404653, 75.4379295410729,
  6.76898432697784, 20.3241143834515, 74.3199198711506,
  4.62053128555435, 18.6060228544865, 83.9066545222218,
  5.502150347246, 18.3315512085137, 83.522710326252,
  4.19489579733071, 19.2869748528168, 83.3107192848557,
  4.92087623242468, 22.2966762421268, 71.4801973059676,
  4.74991983716174, 22.7364458422738, 72.3618869394017,
  5.7959436310297, 22.6131099153094, 71.1139640764884,
  8.59182426714109, 11.0109308738107, 89.1710036921799,
  7.59545039569018, 10.9931867043183, 89.2542157870878,
  8.95078315083514, 10.0823397607021, 89.2651687837632,
  28.1029183981685, 30.5973534704756, 78.6288441536509,
  28.6434425017005, 31.1506335681776, 79.262653925576,
  27.8921153655101, 31.1355856296108, 77.8128366633085,
  21.1722517864606, 30.6580262475656, 89.3061416668884,
  22.0555378171595, 30.1914630219181, 89.3522344477298,
  20.4424325648598, 30.0132717958419, 89.5334203521286,
  13.5050886771529, 2.52193962012582, 79.3624395920829,
  14.4614446719116, 2.28035096568404, 79.198067656114,
  13.3408279149407, 2.58158717725727, 80.3470514805576,
  11.1442872267375, 18.2170700597974, 67.4048732452087,
  10.8566353446432, 18.209231788135, 66.447170286967,
  11.4434158638574, 17.3006020162381, 67.6705956258795,
  3.86891562019796, 1.36091976447153, 66.3795558057917,
  4.2213628094415, 2.26851795156761, 66.6076928470065,
  3.45039222694617, 1.38437641112625, 65.4716527520306,
  27.6800329048492, 29.1944658876954, 73.8907187692247,
  27.5544809015782, 28.2698033636627, 73.5312248038733,
  28.6433242106145, 29.3353207273261, 74.1192571125932,
  13.3474665880024, 2.44635504925951, 85.2015841805407,
  12.6926084425511, 1.77739587083135, 85.5532294946469,
  13.8948887336401, 2.80598615770893, 85.9572259344829,
  12.0298987218974, 30.7040667937021, 82.4030412596161,
  11.4792365664369, 30.0664533403869, 82.9417622214276,
  11.9174102561813, 30.5020157421981, 81.4301477825762,
  25.6393440223669, 10.1136388120303, 71.7648753403184,
  26.2444271760345, 9.70928678970936, 72.450713381836,
  26.1791435324451, 10.6608893736927, 71.1252400444822,
  19.2020304893584, 0.584271301824707, 79.1398326989588,
  18.8501371242971, 0.31031369911765, 78.2447805822947,
  19.7247071428883, -0.169791601290196, 79.5375741400996,
  5.26044049386231, 25.0630002153081, 72.929120099942,
  6.23234708226973, 24.8293364740057, 72.9008563526533,
  5.0010055293428, 25.513808944304, 72.0750328742759,
  14.9230994735149, 15.6899848111935, 67.0954455455822,
  14.952118763252, 16.0226987870045, 68.0380267310103,
  15.6656078352301, 16.107422214357, 66.5715874090384,
  0.291794103783072, 7.76683433664735, 62.881753311353,
  -0.535234402309229, 7.28322643752088, 62.5951398957332,
  0.726174520388152, 8.18582870404209, 62.0844093618798,
  8.00792876486833, 1.66754588584437, 84.232535145515,
  8.38912627376605, 1.69614459007933, 83.3084839708898,
  8.11621328580011, 2.56236038249891, 84.6656419211529,
  16.671269203226, 17.1469701068218, 85.5444260343629,
  17.0973009313939, 16.6264993603081, 86.2844308780076,
  17.2963763450694, 17.8654439054243, 85.2394072448793,
  9.76002614998064, 30.3873535305133, 61.1297979510309,
  9.65435726960497, 30.1545224469866, 62.0965573700509,
  10.5890456469665, 30.9329239230367, 61.0069988450932,
  18.6258960184009, 26.1842056671035, 78.5398434338895,
  18.2576059005781, 27.1133656615135, 78.5718449010764,
  17.8729295446892, 25.5263847436695, 78.5575386919709,
  10.9757433284971, 29.7669250000323, 70.0147657194981,
  10.8867297475693, 30.7599174413035, 70.0924998432058,
  10.8504194111545, 29.4946779588666, 69.0607345542218,
  29.3958268745899, 2.76849177779314, 84.4164610040931,
  29.9892209592828, 3.55827666766394, 84.2611442696979,
  29.1499620358717, 2.35842666934154, 83.5381688614021,
  19.1438618801337, 9.5765085041233, 56.8997787396795,
  18.9929822976155, 9.03014636823785, 57.7236256720947,
  19.2954105475916, 8.96902268498627, 56.1200390517457,
  4.27333017142604, 6.20724627567371, 61.4267086491137,
  4.09655142926324, 5.72085344169202, 60.5710385682001,
  4.796439653161, 7.03790757867042, 61.2360302029726,
  7.48929665021414, 22.2924976639294, 70.2801002956223,
  7.928942891123, 21.7427577899876, 70.9903799967634,
  7.3540369204511, 21.7336237812393, 69.4619531274727,
  17.8728262435789, 29.5311469613459, 75.4110574718923,
  17.3794291314416, 28.712794061016, 75.1163409636065,
  18.639998104998, 29.6989078238188, 74.7919422741551,
  5.21125300257518, 0.945396328498699, 91.1924684215359,
  4.73726940587326, 0.183440477055484, 90.7511490014908,
  5.02937225790673, 0.926594517031301, 92.1756092489886,
  11.991066009293, 4.7659086624407, 64.6446656544156,
  12.1846663545377, 5.31316383148258, 65.4589326169519,
  11.4821807488813, 5.31868881306574, 63.9847642247985,
  12.1651528272799, 2.49880707518845, 82.9098739777031,
  11.7422725086416, 1.66929212883659, 82.5450765135024,
  12.5662366386982, 2.3026842246428, 83.8046742926964,
  29.3843415691297, 11.613193493979, 75.7348556399504,
  29.6515416756604, 12.5764461106108, 75.7622143610831,
  30.0105921881956, 11.077330796064, 76.3011253028345,
  0.581961546736139, 7.06307641136782, 78.5960038211842,
  1.18494731198046, 6.49605762852865, 78.0348462080127,
  0.0342949373277754, 6.47730086765976, 79.1934385852653,
  8.10726799625373, 28.9577876975075, 74.8786132217438,
  7.24312560768946, 28.4848759230091, 74.7065307245884,
  8.8545895192753, 28.4552974742431, 74.4438556838536,
  13.3807195219471, 29.2848090210696, 74.0921591288146,
  14.0976876517407, 28.592474257565, 74.0107387621776,
  13.5485334710034, 29.8446461615307, 74.9035904904605,
  6.93227924959495, 24.8213785700512, 77.415402287656,
  7.9220130148057, 24.775583234203, 77.5507901054843,
  6.65806916688188, 25.773450265315, 77.2798725211244,
  9.95494770956649, 20.8772529967431, 88.5903172875066,
  9.47490918550136, 20.1144838662877, 89.0236142630762,
  9.63417762770699, 21.7391900201646, 88.9829635943006,
  23.1809950583832, 23.0172122248149, 81.8112955668588,
  23.0059526601118, 22.3254802472105, 82.511914600262,
  24.1394802932245, 22.9714967826098, 81.5298419242545,
  0.784508794333807, 8.20388897040949, 60.1244468214135,
  1.71686815228078, 8.48306221318581, 59.8947332428717,
  0.676602664979868, 7.22542605873178, 59.9484735344662,
  20.0387953494842, 5.2826932301587, 69.9678042115717,
  20.4529704398192, 5.92283357322292, 70.614858564565,
  20.1242276362202, 4.35067622277848, 70.3200053222132,
  9.8353507239853, 23.3282088769022, 66.5518319315448,
  10.2465458000522, 23.4058969161068, 67.4600627270934,
  10.5576265032308, 23.2809254134497, 65.8618449948574,
  11.0477468468495, 9.16963137485074, 86.9241132331059,
  11.6058727840007, 9.99934633565858, 86.9158354259827,
  11.6433017457615, 8.36773680309545, 86.9718569046373,
  16.1660456380208, 14.6695329354472, 59.1551604141548,
  15.5314669107615, 13.902558776197, 59.059973871238,
  17.0415722104831, 14.336337422767, 59.5050660746437,
  8.81534613558121, 12.583791227524, 67.9267907652957,
  8.05871559003629, 12.5285244893046, 68.5782934937589,
  8.46922019541229, 12.4347558407051, 67.0005158131255,
  3.30555761737548, 7.16416755912751, 75.8273420507563,
  4.21961201361792, 7.42498843359185, 76.1379495718397,
  2.681313247852, 7.93689278554612, 75.942297222778,
  3.26600594994583, 24.6368606118143, 64.8619551333986,
  4.03490776110268, 24.3909689850366, 64.2717625269721,
  2.93186233540322, 23.8198209261335, 65.3318425634103,
  -0.0378404666901488, 0.632926061566143, 93.7398704373288,
  0.223751516407068, 0.433773204841624, 94.6842791274825,
  0.112773034017498, 1.60306805796635, 93.5497649923116,
  21.0489574060185, 10.9705433110295, 59.9548781277694,
  21.8366691402778, 11.1579433081711, 59.3680293697563,
  20.5398169436844, 11.8171600868394, 60.109849171941,
  29.3913634740894, 23.6973604646915, 80.0410539362086,
  30.2129613150819, 24.2643040412758, 80.1006523308695,
  28.6900856266677, 24.1807451903645, 79.5170800936348,
  7.94834344967438, 15.1202320654585, 85.0403339990417,
  8.94140207164495, 15.217603841523, 84.9743543767636,
  7.67296672825802, 15.1562267144924, 86.0009962948267,
  29.6703503248641, 20.8085989165277, 79.8453712960939,
  29.5376417577684, 21.797732580387, 79.9086408088122,
  30.1347776255707, 20.5887779285478, 78.9874750228756,
  22.5317675150761, 1.90552693161054, 64.6758451948873,
  22.5217271709336, 1.67870648303671, 65.6497300318153,
  23.3416634079427, 1.50386931085063, 64.2483644369539,
  9.95059298403378, 6.29273150054804, 85.6057169383413,
  10.9337846750734, 6.4694885421323, 85.6514449048503,
  9.47591357417973, 7.12286488247659, 85.3132139023426,
  12.4668323689853, 9.88234961420897, 70.3605713485455,
  12.9555935836602, 9.95712127672918, 71.2297788459323,
  13.0243400256511, 10.2760793044223, 69.6297073777523,
  20.1811109360141, 19.5946021036511, 58.2651685274625,
  19.4043847533891, 19.3327401868163, 58.8379902918329,
  20.4691970655752, 18.8105151085257, 57.7154286198428,
  29.0597127140098, 9.6448290524173, 84.9862075901386,
  29.7179198927344, 9.96427976072673, 85.667907344309,
  28.6110131928551, 8.81546212325541, 85.3191028237003,
  8.10446476814507, 21.9622103148214, 62.3272216112453,
  7.81519184594862, 22.1687241339962, 63.2619264946036,
  9.03491965327378, 21.5960081901648, 62.3394572410677,
  2.98832347887578, 2.23485420525403, 89.2623242757506,
  3.53892059815382, 1.45726993027708, 89.5659778737061,
  2.95679898491779, 2.92394772397752, 89.9863106904947,
  29.9277174237296, 23.1724759286993, 71.0744162780346,
  30.2716344341012, 23.9586132649338, 70.5608900581051,
  30.6542468488594, 22.8132338031068, 71.6601637403598,
  28.6280370592425, 7.35633051010593, 62.2474398052178,
  28.4315712651332, 7.95807659044429, 61.4732932773935,
  27.7697180600113, 7.06941454509058, 62.6728428195208,
  13.9620944762963, 3.011749703545, 69.993275408273,
  14.4199613909609, 2.75505566196754, 69.142119689574,
  13.2998458322086, 3.73816993957224, 69.8095898778301,
  9.31806872167112, 29.5084105192097, 93.287436489049,
  9.90988041641716, 29.0489653011951, 92.6251155626052,
  9.86859659548197, 29.8364315156056, 94.0551091315736,
  4.46601884347906, 2.03807838154433, 75.2403113463103,
  4.34624213781106, 1.38336937266653, 75.9866421405789,
  3.61928842858598, 2.0997470602753, 74.7118753723659,
  25.1730872551366, 23.5613488174852, 88.4820506113807,
  25.001864924448, 22.7221568530258, 87.9658725798252,
  24.9059462003518, 23.4261979612435, 89.4361836749025,
  23.8074077349457, 16.9270377816096, 80.1969718565488,
  24.7061616031011, 17.0721943113139, 79.7832436047218,
  23.5262666236789, 15.977376043752, 80.058760933663,
  5.28568766230325, 3.7698483408189, 80.3529629207053,
  5.29811320506512, 2.79232218785873, 80.1425152403523,
  5.52236778210638, 3.90678379493178, 81.3148523126298,
  15.122537819238, 5.17795245457702, 89.6612397733439,
  15.0062333483045, 4.26666970050085, 90.0562549783224,
  16.0967849269797, 5.39791643742201, 89.6116573237464,
  7.39898563805368, 14.4814668444475, 80.6596793604438,
  7.30612631782125, 13.7072458119968, 80.0336131182961,
  8.0715556721082, 15.1257531975434, 80.2956125471989,
  7.57556362995432, 0.389275656756873, 86.4582925272668,
  7.69555196220103, 0.836254758583539, 85.5718318780246,
  7.37423271749149, 1.07829851056348, 87.1545061228099,
  18.0544956481205, 10.6400591915063, 71.8701079455886,
  17.887714094841, 11.0314673801011, 70.9651308500846,
  17.8080292029722, 9.67092285172789, 71.8647184802362,
  29.4274422585045, 8.73722932320605, 91.3338705098411,
  28.8051409211389, 9.48384155989807, 91.5690538713588,
  29.0615105766283, 7.87524194304441, 91.684686359884,
  28.7395218859489, 20.5533865610046, 70.7882184167185,
  29.0853102461392, 21.4503570622952, 70.5127654628928,
  27.7814940663738, 20.635432531832, 71.0629021541171,
  0.689501388503436, 20.7674130154485, 63.6865720007293,
  0.130339535322376, 20.1965394561621, 64.2877719685062,
  0.101628712717085, 21.410984302382, 63.1964478167734,
  12.3649915376852, 1.1192438722163, 77.1846773830682,
  12.559981348388, 1.67746610571841, 77.9911306748006,
  12.619997296896, 1.62426505038821, 76.3601013269235,
  15.6452353778094, 16.703385365906, 83.0602459803566,
  15.8863534309762, 16.7806294526638, 84.027662868517,
  16.0758705493067, 17.4471186729404, 82.5489592534829,
  7.25315517409302, 28.8175873142547, 90.5705549784973,
  8.24280311156481, 28.9303498781185, 90.48177680523,
  7.04812147264512, 28.3282241543549, 91.4181898521331,
  28.8820167838508, 12.5548394420751, 66.1214708851009,
  28.7586199874936, 12.0360936281754, 65.2754945194676,
  29.6896030120297, 13.1388760694733, 66.0395825348105,
  7.59323645390827, 21.1447804632024, 84.8515192518156,
  8.06745705096801, 20.2818856846198, 85.0262402477468,
  8.24063258764038, 21.9028445608614, 84.930367649828,
  1.48250793053232, 17.2170796134708, 78.5961181419983,
  2.33018035730086, 16.9264066020209, 79.0399206400884,
  1.62601277258911, 18.100094778935, 78.1492506248676,
  9.77730545719679, 13.425905613507, 59.3153629737073,
  9.3144618341313, 12.9381369666984, 60.0555369585096,
  9.94822951775531, 14.3708031030533, 59.594564871572,
  7.82047830918158, 15.1892727859708, 69.4027421988183,
  7.74156637495836, 14.230803675044, 69.6768039984845,
  7.20416811035584, 15.3685382250658, 68.6359138991517,
  18.6528578433705, 24.4149516262501, 66.098310663972,
  18.4633170304582, 23.4418680979587, 65.9672277619274,
  19.0769607202219, 24.7861818837692, 65.2722810968567,
  25.0058511942293, 30.71658628737, 81.0409108987652,
  25.456387367088, 29.8349919905012, 80.9001676833897,
  25.6930494401367, 31.4127358231947, 81.2485991136278,
  24.245881840613, 26.1050023186745, 87.4911819398584,
  25.1099656257565, 26.511483715826, 87.1943114529087,
  24.4114660333863, 25.1772989614378, 87.8257687837052,
  14.711690823284, 26.3344098320859, 86.5930510992979,
  14.8085649284444, 27.2862070379958, 86.8840794253618,
  14.7795885227632, 25.7337042260636, 87.3896329703563,
  23.3259134717076, 16.0397581254937, 84.2468822494121,
  23.4072655655877, 15.0430761355953, 84.2494990859549,
  23.3876753388724, 16.3817154654893, 85.1845659110952,
  17.3983216864351, 12.2192720983753, 91.4921939181804,
  17.9705154816303, 11.4006498199464, 91.4426780015478,
  17.9079425356102, 13.0040229606662, 91.139415412288,
  5.58082442445091, 28.1807732273842, 79.3054016389849,
  6.57309619016128, 28.260989945729, 79.4000695906476,
  5.21572688309034, 27.6438716085955, 80.0659543571015,
  16.3069341017689, 12.4308674355811, 82.9989297126678,
  16.9590333884366, 12.3994471644149, 83.7564119150246,
  16.4580194141792, 13.2616664836528, 82.4632561459342,
  2.72966788221601, 9.4589485060478, 66.5392291245318,
  2.73849212883974, 8.46005860046256, 66.4929572195415,
  2.59495919388631, 9.74756255049742, 67.4871507999011,
  30.8532973713659, 2.85676830685592, 61.8233243111881,
  31.5542419210193, 2.16168935740881, 61.9831429344671,
  29.9582774140213, 2.41685408476504, 61.7497393048556,
  5.4592883904622, 17.8038936571538, 86.7585206876954,
  5.82957207145144, 16.8858137432482, 86.9000101476426,
  4.51843228196318, 17.7363458135715, 86.4265160613308,
  24.0479273383553, 29.4047636284489, 88.8753509930487,
  24.9724052122012, 29.0385253770888, 88.7694727421662,
  23.3808040623914, 28.7041340469507, 88.6222408901354,
  14.7447434238252, 3.62099329300326, 63.7620712470911,
  15.5464173214798, 4.16493721177897, 64.0099501994976,
  13.9377206067167, 3.98604393804328, 64.2262395347004,
  28.5230983825991, 9.07537079860653, 72.3068689230725,
  29.4893196636844, 8.82312902643993, 72.3596943369575,
  28.4377399884131, 9.98460042869071, 71.899419019012,
  7.43885454486813, 22.4119990589467, 76.3529045290498,
  6.86011942579379, 23.1412126817702, 76.718025268311,
  8.30587147673613, 22.3936507411996, 76.8508452675821,
  5.3646161880913, 9.22666788939009, 72.3973517829415,
  4.88903611167012, 9.85218566715414, 73.015858937801,
  6.24183297566704, 9.62528229612438, 72.1297751353447,
  26.1316498261853, 27.5071765293641, 61.0436323462137,
  25.7458945289489, 26.8369893068402, 60.4095645758454,
  27.1189808099055, 27.3666141850883, 61.1172513380428,
  18.0343719707574, 0.727113689205625, 85.0210621142551,
  18.7011825903021, 0.315453800509021, 85.6422703995353,
  18.0912365719279, 1.72352769855046, 85.0837162371448,
  8.17667981241079, 2.27340423699811, 61.6618656423532,
  8.85901983195673, 2.77170405225366, 61.1269736982726,
  7.44873813056388, 2.90000810525785, 61.9401972792755,
  28.1261705467085, 24.4456739493738, 92.6883023100813,
  27.7286373811125, 25.0235585666526, 93.4010552485977,
  28.8732803069778, 24.9361303559093, 92.2396604491291,
  28.73038201813, 3.13986589435477, 73.4178135557743,
  27.7770236490849, 3.05045228056581, 73.7061068540676,
  29.1806572188047, 2.2487573985858, 73.4741863544074,
  27.1145779388047, 13.991132613191, 84.6727453088957,
  27.6993716652813, 13.9134895165471, 85.4802029529966,
  26.173067947803, 14.1690967128687, 84.9589056067532,
  3.66437043811507, 20.7762720912386, 63.286000464599,
  2.69338810802502, 20.5384675524375, 63.2606565111099,
  4.21106294517302, 19.969845979572, 63.0606025294955,
  25.4440087806173, 4.12736270576344, 69.9162536890468,
  26.419924166482, 4.34496800858658, 69.9316514751133,
  25.026003388491, 4.40904133276463, 70.779925295182,
  14.1599140676016, 11.0376355461445, 68.4019696054802,
  14.9509413901865, 10.5818728068164, 67.9938567529943,
  13.5611991170027, 11.3788029069694, 67.677300550092,
  1.76852145440544, 4.22299612129122, 66.2408722712797,
  2.47045660110693, 4.79983006144016, 66.6586636729593,
  2.15221321727228, 3.75465154578326, 65.4449866075689,
  2.94885978668948, 25.0284636624141, 80.198478771625,
  3.38438551403489, 25.7103311308741, 80.7861641434663,
  3.54088179133058, 24.8359512714064, 79.4158876105906,
  21.2807826048008, 15.4488076960054, 68.0145845546848,
  21.4099693159844, 14.4801966080567, 67.8022090524338,
  21.4921647855173, 15.9983670096974, 67.2063134773785,
  20.4746397386713, 0.3407782210638, 86.6672967306514,
  20.828293842272, 1.21607274928478, 86.3374660712627,
  20.8736024961979, 0.135509230516283, 87.5609931889786,
  29.5166371483591, 30.7082963427909, 89.1851545043009,
  29.5698400236289, 30.1792512635323, 88.3382302112408,
  28.5594409742301, 30.8059290634289, 89.4576308080295,
  2.32387793154697, 3.40575590401911, 84.8520919828045,
  2.72082158393952, 2.77381716550959, 85.5177414157617,
  2.08152744003094, 2.90544335277974, 84.0208558007634,
  25.1109274954196, 8.89299037459255, 67.5506825547687,
  25.6212578759944, 9.53492299215042, 66.9784191388686,
  24.1879997821402, 8.77948932958772, 67.1828212373626,
  2.68893644503877, 15.92407257331, 72.6621630825029,
  2.452083455626, 16.2270973096541, 73.5852430739283,
  3.25123690108435, 16.6207201016161, 72.2166292247144,
  8.65754813276055, 21.6192852964099, 79.2582679294864,
  8.90944651758536, 21.440252604904, 78.3072187724525,
  7.73065904990819, 21.2837325896441, 79.4264375137495,
  14.6122531580311, 20.9081091951965, 67.7776711611813,
  15.2186594083337, 21.1187082251875, 68.5444302551352,
  13.6834439330778, 20.7611709520912, 68.1178513727676,
  12.2747024413103, 26.9186436216615, 69.2570452491072,
  13.1816011618714, 27.3232475053867, 69.1394424943817,
  11.7993829382592, 27.3782328399919, 70.0072779599468,
  10.428340885404, 28.709868085807, 88.2907889404045,
  10.4588343443186, 27.73330959852, 88.5038703095365,
  11.3581296119342, 29.0490408624239, 88.1477688312609,
  6.02830855854286, 8.02527133038081, 67.4843212031003,
  7.01696788508115, 7.87628386040571, 67.465467295301,
  5.77256191695743, 8.456051751219, 68.3497817073061,
  23.2863187891168, 0.154978369373597, 72.7662844820051,
  23.3166701776687, 0.791520809612252, 73.5369287027633,
  23.9343271650208, 0.450332700248941, 72.0642510326657,
  10.2535747402433, 24.7411674876953, 74.4267539417064,
  10.060482324929, 25.6723322887536, 74.1174847508416,
  11.0455624649093, 24.3831558620061, 73.9322004867091,
  15.0003084117448, 5.79482151885779, 84.5710198684869,
  14.1131127910184, 5.90433040002181, 84.122810391222,
  15.6542214828447, 6.44153125310027, 84.1783823574404,
  21.5671683112252, 17.6484880816274, 56.6993739350507,
  21.7774057498752, 18.0164982333413, 55.7936318373069,
  22.3897996594974, 17.2360984137891, 57.0907975249121,
  5.93509303096998, 8.45562714794059, 76.7322154271704,
  6.78426085452096, 8.52023991939123, 77.2563711265681,
  5.23069303562215, 9.01559532094688, 77.1683992092783,
  2.50035189190577, 6.35680043921269, 63.6647273518346,
  3.09293181620486, 6.41828257075343, 62.8615654871903,
  1.67445550381305, 6.89953179069079, 63.5119600900992,
  18.196298926855, 5.53641995357108, 75.1237573284473,
  19.0095738498522, 5.19549916796431, 75.5953046935817,
  18.4713547436188, 6.169322625066, 74.4000318928856,
  24.0759418455356, 15.381018689867, 69.214564326612,
  24.0857292210688, 14.9763671789265, 68.3001457342956,
  24.1818345916262, 16.3727007955911, 69.1413978895515,
  30.0312322828584, 22.2152900503804, 88.4729014479824,
  30.5275505368726, 22.4185335795536, 87.6288870769071,
  30.3564143173867, 22.8155464994779, 89.2036194782354,
  25.5965820135313, 25.3899908071229, 59.4303470402221,
  24.8565714043934, 24.7536879511243, 59.6482988096836,
  26.4292115321398, 24.8753990099237, 59.225595075648,
  30.305882770639, 5.33524288248571, 80.8588817041526,
  30.6343627648663, 5.13102200211044, 81.7810501949455,
  29.7025698815818, 6.13218630011374, 80.8887940259761,
  30.1991211343334, 5.29754080454636, 87.9138082152922,
  31.1417772233687, 5.56977855742575, 88.1069043149726,
  30.1418154607513, 4.29999215361856, 87.8736491713865,
  25.3695970716526, 5.80396330591518, 91.8249377065342,
  26.3649282481477, 5.70759454319694, 91.8195608422817,
  24.9748153839923, 5.14958399541236, 92.469868041589,
  6.7100483431821, 17.8512564760367, 76.6332594518353,
  6.6993523199706, 18.232239467883, 77.557779627392,
  5.82143012101372, 17.4389703331347, 76.4323171924638,
  18.553759203447, 16.4489944125917, 61.9550836659496,
  18.7564740604436, 16.6018194512586, 62.9223226200397,
  18.5110692125909, 15.4663327554456, 61.7746574143799,
  13.8947293537474, 9.7972379666396, 61.4422644030235,
  14.1663933785096, 10.4658723557952, 60.7500746087557,
  14.3839352434649, 8.93903003790173, 61.2868399888628,
  30.4399107608698, 9.0189189082872, 65.3782998374577,
  30.3821190276751, 8.3215647627986, 66.0926928044893,
  31.0663317462485, 8.71130119190286, 64.6620819309212,
  31.2325245219715, 5.4928356820712, 73.4703629559155,
  30.998490793803, 4.54577532348947, 73.2505792183856,
  30.4781778647989, 5.91444917377288, 73.9735559451629,
  24.7400286244241, 12.7558068536167, 67.0822790039958,
  24.6401731101226, 12.842374014976, 66.0910499674771,
  25.5608703251891, 12.2235276206954, 67.289396652896,
  23.6935870739514, 8.53532510762671, 70.3310732687221,
  23.9056602624654, 8.57718320900214, 69.3547163349818,
  24.4247207229492, 8.97790354520031, 70.8502725694711,
  6.9519537977036, 16.319926842258, 66.9265044589102,
  6.92305298069202, 17.2936698911574, 67.1523123805961,
  6.14112786931241, 15.8674396889664, 67.2977411623147,
  2.15131496397892, 24.7178207459715, 72.3859489092544,
  2.09596231269408, 23.7212961335655, 72.3237011714252,
  3.06460279755667, 24.9822461190308, 72.6957626518826,
  26.8301604041068, 7.14763707529052, 87.8439784681392,
  26.7991530722094, 8.13452117726767, 87.6855539920209,
  25.9763938147817, 6.85181729017648, 88.2724329764445,
  2.04456335100659, 22.18854075295, 66.1496471910135,
  1.19605027209715, 22.2536594751277, 66.6747996516776,
  1.89039122915135, 21.6292496259638, 65.3351385095883,
  26.2817614043243, 17.8217109830327, 59.1138322628246,
  25.5535721210755, 17.4472308574166, 58.5398069991993,
  27.168064522718, 17.502030087486, 58.7787637514002,
  2.76204698049934, 27.7310889299368, 75.5221034262273,
  2.11740215080536, 27.0178392688311, 75.246952623064,
  2.83773604123215, 28.4113036661514, 74.7930087281792,
  21.143761647302, 13.4022909424351, 88.2852849727859,
  20.8605878104257, 13.1279153564864, 87.366301503977,
  21.6744487566088, 14.2481783558475, 88.2319400963124,
  22.6258153479058, 2.51862992040298, 74.2620251745708,
  21.6684040785237, 2.42141694398637, 74.53389517747,
  22.6736348025264, 2.92551548356631, 73.3497985370245,
  30.5214985415744, 17.8386088928469, 67.3351949025479,
  31.1929492639045, 18.4048982760106, 67.8131805320374,
  30.5080195301607, 16.9242903160713, 67.739966265683,
  4.99491202736656, 28.2967741220245, 94.6657279513058,
  4.75728721154017, 27.7166577028671, 95.4448296052171,
  4.42525308412523, 28.0513142791682, 93.8813567675349,
  16.8630372790225, 28.4650520179178, 86.0385241865174,
  16.2089987290265, 29.2199687224298, 85.9902091332958,
  17.7903612656537, 28.8317007464459, 86.1136170203105,
  23.2830412081009, 18.6044083883889, 71.3973152810256,
  24.1371502046246, 18.1378911670426, 71.6272272299204,
  22.5096753537175, 18.0747226011317, 71.7456516444039,
  23.7608675145372, 28.1525767209084, 72.3712284355987,
  24.2026287458098, 27.4938281271826, 72.9802418219941,
  23.676674772411, 29.0332060734873, 72.8374939453137,
  29.5232722004008, 18.5702182997006, 85.1554284814496,
  30.0667633840063, 19.3123626095384, 84.7632051308974,
  30.1303819239985, 17.83247752719, 85.450651001066,
  11.8569003335178, 6.14730723811089, 79.3151624457198,
  12.3465171125188, 5.69198612118204, 80.058773964054,
  10.9683191067011, 5.70804278352293, 79.1829877799002,
  9.7435515274547, 4.18659169945868, 87.3374398052759,
  9.92294098243277, 5.00294770841235, 86.7884568455332,
  10.5776517651025, 3.91955523146146, 87.820107722498,
  3.50749728461687, 23.8691493753477, 77.3348123419576,
  2.52115761819775, 23.7614882348806, 77.4594844771022,
  3.71725628853243, 24.8292003823831, 77.1496010459556,
  19.6614120699201, 14.1244126108691, 71.6857166982356,
  19.8543940147431, 14.0711916827294, 72.6654745773977,
  18.6720430577595, 14.1413611720628, 71.5412808853292,
  13.9958384269121, 17.6555946516937, 86.1423354388027,
  14.9929482782341, 17.5814642014637, 86.1257035193333,
  13.7198715666254, 18.5299319654608, 85.7431155072136,
  22.4335932568793, 29.3292118319297, 77.8700300286978,
  23.3249908150417, 28.9613114476371, 78.1347179591734,
  21.7997352805453, 29.2532630125778, 78.6397415608167,
  21.3769352864907, 19.3650019955049, 67.3481161593568,
  20.4655566348367, 19.1613084047866, 67.7057442824255,
  21.8399829604371, 20.0054496709004, 67.9608262267895,
  13.1597861355372, 29.5511555526902, 85.183763457925,
  12.5412699665443, 29.1315833960281, 84.5193863405825,
  13.9072706705373, 30.0077390949276, 84.7012716560325,
  23.8067198938895, 12.4238624886111, 56.564021615084,
  23.3888287974451, 13.3230923990888, 56.4345897812304,
  24.4817651480251, 12.2632251870969, 55.8439455342207,
  19.9105904492205, 16.5616418865034, 84.8198849102012,
  19.4464123021372, 16.7513053233957, 85.6850822451927,
  20.7632566746184, 17.0824081688642, 84.7778993505197,
  23.8203710687765, 11.035187418071, 58.8510007241758,
  24.0943677845123, 11.2592707561742, 57.9157400881227,
  24.5302332609676, 10.4780246596846, 59.28188972237,
  30.9377636249076, 10.4767595558176, 73.6439968474292,
  30.3948192683545, 11.0107767297725, 74.2920995272635,
  31.3330236517644, 9.68637526131514, 74.1120376342982,
  23.5740983816759, 0.930231964113279, 78.8824118196002,
  23.0506561925242, 0.199564403915346, 78.4440818171015,
  24.0638375821727, 0.561616050488205, 79.6725243582421,
  17.6119134874623, 18.7319717852456, 70.9745277382015,
  16.766471064241, 18.5796287689463, 71.4864053743632,
  17.41912445785, 18.6952952159299, 69.9939731913637,
  0.189835893000315, 2.74329052975538, 89.621800204877,
  -0.477119021620813, 2.72102024877437, 88.8770350227909,
  1.10068471805036, 2.54535975755131, 89.2596154076813,
  19.3152426675776, 2.37574959428349, 66.2814044244304,
  19.8639636986801, 3.19574073567957, 66.4442533054758,
  18.9657521500587, 2.38915497531186, 65.3445604278526,
  3.42202965633876, 3.71407742453742, 71.5263164289166,
  3.21745135071987, 4.22356791682264, 72.3621197282288,
  3.23294707986681, 4.28936414941065, 70.7305193671858,
  25.501967277316, 11.7169303724939, 88.1203278813425,
  26.1203032640474, 12.3454450108942, 88.5921646718002,
  26.0071999539982, 10.9014160535313, 87.8380579077719,
  4.7732704796741, 19.9606743755539, 70.1537274015795,
  4.74876452766899, 20.7858801769643, 70.7180277149189,
  4.40343204895128, 20.1654569049281, 69.2474803873369,
  16.3095334647405, 10.1246800465013, 66.8022717277358,
  17.0875682333365, 9.50227199727737, 66.8875367212384,
  16.1780447139446, 10.3641038204632, 65.8403013722279,
  13.1341818993197, 29.1494645544948, 87.9568492431883,
  13.9699916373448, 29.5042095767341, 88.375869589972,
  13.256246835597, 29.0926262589878, 86.9659559293066,
  20.5806834557133, 26.6788024220834, 80.3572126311342,
  20.1707722068832, 26.5653481814031, 79.4521706965509,
  20.0300328176592, 26.1927758179999, 81.0358598258781,
  7.43243240018357, 24.3909808732046, 87.4324013048286,
  7.48772813798619, 23.8917210333255, 88.2970873713665,
  6.47636600807863, 24.458842318838, 87.1472138610587,
  7.67591314520725, 23.4329672426045, 73.8009464433554,
  7.08400854740001, 22.9165122666437, 74.4197543334958,
  8.38973022260552, 23.8930067813596, 74.3289888685417,
  13.2332320385836, 27.2959784557804, 90.0159433366082,
  12.8668897004512, 27.766878988632, 89.2134185834375,
  13.4894224606498, 26.3621182308569, 89.766400659001,
  6.64697154393532, 29.855871188659, 71.7147206696559,
  6.92408588910294, 30.6416721551783, 72.2676442454959,
  7.29728655468123, 29.108102045241, 71.8486299484621,
  17.3797728561993, 4.97316558651529, 69.1476537636793,
  17.0621977145606, 4.0657768723897, 69.4229567801732,
  18.3308040854764, 5.09399977686398, 69.4321510385035,
  18.9214485132687, 16.1136933036576, 82.1099482291041,
  18.7963486678191, 16.3436976623895, 83.0750637784726,
  19.8975525584934, 16.1066446267706, 81.8927588899317,
  27.9667683672342, 10.5833787097901, 56.1326439729548,
  28.6590289759068, 9.94717515330517, 56.4732614774905,
  27.4312813990626, 10.9356227112153, 56.9002232003824,
  12.4431608756949, 1.83512603572148, 73.5608759792347,
  11.9638457030925, 2.66519734453506, 73.2758521423408,
  11.7777406524089, 1.154740620597, 73.8679453742058,
  18.8503765337067, 29.067899600231, 90.1081427687406,
  18.2397363896807, 28.9439529100329, 90.8902909851886,
  18.5657400202798, 28.463595737865, 89.3639661115188,
  26.5076933541098, 12.172527402159, 57.779944996599,
  26.9662004674662, 13.0355735314916, 57.9918945322097,
  25.5507838897105, 12.3509279374921, 57.5508216107655,
  11.610641796334, 12.5915433898921, 71.9291846065818,
  12.5142159920155, 12.192879600782, 71.7722742622734,
  11.664387726802, 13.5858266397381, 71.8369230542767,
  7.06040965921238, 29.6773324857882, 63.5420488889591,
  7.76514107036566, 29.0592249135705, 63.8903255997814,
  6.79027774440542, 29.3907258889539, 62.6228724057668,
  9.23549853737475, 18.4477389727038, 81.4061686635018,
  9.40516889011205, 17.5732665025671, 80.9517350925863,
  9.8556226193257, 19.1405327536646, 81.0380886449643,
  3.81547654842287, 14.3208320595736, 87.6411060961733,
  3.38212555678771, 13.5044856391981, 88.0229246918298,
  3.20349497580828, 14.7405071895495, 86.9707693598535,
  13.3649218089162, 11.0705633254546, 82.3867574253914,
  13.4421366793363, 11.1717972640433, 81.3948957649448,
  14.1682552444583, 11.4722960247893, 82.8263779772603,
  15.3359628175238, 6.46337827028928, 69.6903327405788,
  16.1567892289721, 5.94670183717813, 69.4468384578196,
  15.5998564079645, 7.30989437746984, 70.1526861262138,
  0.442440316303067, 28.6399299729331, 79.4991727468709,
  0.236440217196698, 29.5653713968253, 79.8171698067827,
  1.07443470336338, 28.6862272050587, 78.7255839277804,
  26.159254706666, 15.1987347382183, 80.0180458390261,
  26.712077812867, 15.113871887466, 80.8470120083072,
  26.5606466684069, 15.891738057845, 79.419187849152,
  2.24620376147696, 5.86288384319089, 86.4864881387225,
  1.63442707495198, 6.47116200409821, 85.9807936016868,
  2.43842083029863, 5.0505028994514, 85.9359522173672,
  20.1466321770387, 4.67645331067979, 76.94278478542,
  21.1133678770772, 4.68787181777384, 76.6872623715955,
  20.060189809852, 4.82987206934428, 77.9271578862538,
  17.1981910558114, 15.5007902813187, 73.6584019364839,
  17.2779036964972, 16.2299494813552, 74.338087713823,
  17.9441485677748, 14.846450589426, 73.7824461139341,
  16.7353435885399, 7.83740547158428, 72.2705913241583,
  17.5793030996187, 7.3284861059012, 72.4401006834644,
  15.9765567495493, 7.39255060463232, 72.7463503811651,
  3.55662393844962, 22.0397997884147, 60.738267800079,
  3.5779118151575, 21.6654165413498, 61.6652974709215,
  2.94604512461164, 22.8313316506218, 60.7123675451926,
  15.3257869194361, 27.1384681235764, 74.3396112161316,
  16.0870036244407, 26.514965314513, 74.5179181849016,
  15.1512905876005, 27.1787090086952, 73.3557760158359,
  22.0101591727605, 27.5137989514253, 88.1533003808351,
  21.4901501793311, 27.7271655304428, 87.3262179486006,
  22.7330614363278, 26.8589455776448, 87.9328930847274,
  1.93378306437047, 9.60751852364062, 75.9672169637594,
  2.6435732524841, 9.91919437625013, 76.5989257983959,
  1.03866440567241, 9.68754747974811, 76.4058032757151,
  3.65497525263551, 26.4969779533521, 87.6412723522137,
  3.382808478361, 27.3366353201476, 87.1712715507602,
  3.36295438455691, 26.5401309290869, 88.5967102797066,
  26.774454442399, 11.8056562257112, 78.6367768131444,
  26.1051480124567, 12.2848452773274, 79.2045855447161,
  27.6120151859488, 12.348887229247, 78.5785352673052,
  1.05821113945219, 13.9735758869583, 71.6548154559252,
  1.67058185060986, 14.6914249881082, 71.9860174790087,
  1.45007448937422, 13.0779059166377, 71.8650972175063,
  20.777874365195, 28.7844512794564, 83.2400446485236,
  19.8514243330077, 28.4215889856886, 83.139938237032,
  21.4376495203894, 28.0354912824055, 83.1787611482503,
  16.8266898786735, 9.10845105334009, 85.373692265235,
  17.2846037235966, 8.82919593413311, 84.5296949376181,
  16.9844190321697, 10.083208750695, 85.5317079150448,
  8.95143945804804, 21.3986405802912, 72.5317038629449,
  8.68970087579585, 20.7746992133693, 73.2680394421506,
  8.51010892774715, 22.2847898005648, 72.6730082239279,
  10.3300188871356, 13.8051781114987, 79.1123443729772,
  10.6457422208979, 13.4372665922058, 78.2377245181319,
  9.95036806392505, 13.0652636141154, 79.6676747152038,
  18.6083085367781, 19.717876493267, 78.507211283374,
  18.134220765153, 20.5021281221406, 78.9074489220399,
  19.5695571740022, 19.9498967999836, 78.3583232895472,
  11.0370370513222, 20.1079797653206, 86.1356601219668,
  10.8606771006749, 20.4419510651086, 87.0615976677687,
  12.021106954637, 19.9847240567024, 86.00754120969,
  23.7416842980542, 0.899640375285258, 85.1725309954042,
  24.2303908088968, 0.616002463562865, 85.9975858307295,
  23.2492815844137, 1.75111555679923, 85.3528905886208,
  10.174738574833, 18.2087108390013, 77.4482859581379,
  9.97398622132974, 19.1882341235161, 77.4330338220164,
  10.1417436984338, 17.8471272309006, 76.5165302860412,
  9.80827106021833, 29.350390722081, 67.3880421593652,
  10.0679957947499, 29.9046532709694, 66.5972602114351,
  9.47248399173566, 28.4615377998616, 67.0762930177437,
  3.71804298410573, 20.6507878469788, 58.2172123658989,
  4.65435448670231, 20.983137979981, 58.1037920890576,
  3.32757815930958, 21.0335634814112, 59.0544817576013,
  14.4538642314103, 5.99538788660989, 77.9953573099948,
  14.5734948000999, 5.22406340012668, 77.370259666753,
  13.4785096064473, 6.18542282827933, 78.1074736625395,
  21.7767278107448, 29.5369754000092, 75.0448069092347,
  21.8337626098628, 29.4041517990642, 76.0343042173268,
  22.6982857910588, 29.5523651662963, 74.6568712908478,
  27.7535202864217, 24.5695214244204, 66.694862853155,
  27.3060623319066, 24.6092619408198, 65.8014413007523,
  27.1190295829544, 24.8864159798612, 67.3998446883433,
  5.55969603297666, 22.2734860513142, 67.0631094107268,
  5.8048419936795, 23.2320174821515, 67.2084399100996,
  4.57844069926514, 22.153779825699, 67.2141338776574,
  29.0592844522054, 17.5723362117829, 61.9345468776641,
  29.367240096913, 18.4966476885976, 61.7091325597484,
  29.2582266495719, 16.9590062906839, 61.1701854382968,
  25.3283593738395, 5.13019810524798, 79.8141270238174,
  24.8637946247111, 5.86456674267106, 80.3089828596288,
  26.1069429098117, 5.5069795126359, 79.3122869610885,
  12.9484663483169, 14.4289665713657, 58.6634854439348,
  13.2956262443377, 15.2550298578607, 58.2195266020361,
  12.0024074031769, 14.5777135690743, 58.9513166496667,
  22.1683385604888, 23.5899524105207, 85.9022354939802,
  22.3345472521972, 24.4422487839375, 85.4062863406779,
  22.8308515325849, 23.5025325470527, 86.6461671637428,
  20.612378916178, 2.42169435289804, 81.0647645506634,
  19.9866360179188, 1.78889198366462, 80.6086867209339,
  21.3782347858711, 1.9102594381738, 81.4545069205152,
  28.3766119007383, 1.88976492217655, 62.5121204756703,
  28.0925602073359, 0.996753773040229, 62.1630564084943,
  27.7489669470201, 2.59312349436839, 62.1784312025488,
  8.80540223397622, 23.2499090787418, 58.7621505263402,
  7.91428196526411, 22.7966572980584, 58.7405290093312,
  8.82517901042414, 23.9106850852951, 59.5124730891602,
  13.4183558119463, 19.9021801745209, 84.4553800075655,
  13.9178716134568, 20.7178456985894, 84.7472253722493,
  13.8106807832869, 19.5585229848583, 83.6021620677309,
  19.1471359229786, 8.8358645199509, 59.4925562332624,
  19.5591553923608, 9.67610736491499, 59.845021718575,
  19.2007652072916, 8.12056637661278, 60.1893147753708,
  28.5938918073479, 15.2754494759904, 90.6668528465494,
  28.1074392977553, 15.889784696498, 91.2881065731015,
  29.0592075085985, 15.8126807735125, 89.9633872602324,
  3.32209984402253, 12.3000229675929, 83.6039813133058,
  3.86578199424344, 11.8117912841921, 82.9213104241837,
  3.86340932358902, 13.0476890414107, 83.988662336224,
  16.1732766742255, 21.7039765861005, 69.9014932744323,
  15.9255146478549, 21.4441541004492, 70.8348240058661,
  17.0619833603974, 22.1624084002384, 69.9078727524303,
  28.8971531616273, 7.09508245146267, 86.243085771457,
  28.0546717058219, 6.94324135696306, 86.759969973813,
  29.6612350466196, 6.65421638529143, 86.714059215215,
  12.8276809443575, 19.1055871514761, 73.7489973869318,
  12.1544653391768, 19.2938398199513, 73.0339157959556,
  13.1386280093201, 18.158202462828, 73.673009397709,
  13.4563869096847, 6.01082517491964, 66.8861413694929,
  14.1607703730613, 6.65010265857554, 67.1946348627988,
  12.8845607577505, 5.74493360169509, 67.6622319075438,
  9.59913142439363, 7.39454229978442, 73.0594233385514,
  8.80804852835072, 7.1596411860048, 73.6242324375694,
  9.37336856353634, 8.17631172200159, 72.4781594560129,
  27.3010985679879, 7.14327197606013, 67.8081746432441,
  27.9809938081866, 7.72070991151228, 68.2601789497014,
  26.4642229826874, 7.66946077768514, 67.6572952219425,
  21.1617208553156, 20.7115942098945, 77.7638532466777,
  22.0690223360712, 20.30437519965, 77.6590834957269,
  21.2437013992001, 21.7080547038704, 77.7824455668578,
  24.8390847257496, 27.2926010958527, 65.8081015570759,
  25.5387388450092, 27.7774107491697, 66.3329288748232,
  23.9791121394202, 27.8012578803956, 65.8495192622315,
  5.08242361450639, 10.8895549397249, 81.9816098531237,
  5.41267901637601, 10.1864535656951, 81.3518640096493,
  5.79877017928441, 11.5726200836312, 82.1239812277431,
  3.09466374447172, 11.7753727358095, 88.5499377851969,
  2.78315969048681, 11.1561826623098, 87.8291265219453,
  2.57407233958549, 11.6023254968778, 89.3860234520138,
  16.8506131538576, 14.8102752258921, 70.7999347515423,
  16.7195815975694, 15.2153188634763, 71.7047940681818,
  17.4590403166841, 15.3914357224008, 70.2595007918092,
  21.5426866135491, 13.789043175066, 80.7221201662768,
  21.5668329443248, 14.2713995127558, 79.8464779344261,
  20.5936248648087, 13.5923771650656, 80.9682995268827,
  11.1875177413896, 0.0723567812092112, 91.4201172427996,
  10.3883313239861, -0.372707927022534, 91.8241203068032,
  10.9374807686399, 0.468231788415225, 90.5365084544052,
  22.6519901180271, 0.716386570172025, 82.3358449411659,
  22.6911682418733, 0.745706616082489, 83.3346469283083,
  23.1387818650658, -0.0927712241222286, 82.0067591484797,
  18.4793484902567, 6.73603724592269, 86.7284970373573,
  18.3699649217632, 6.27330119147175, 85.8487751615041,
  17.8817189667465, 7.53717768535175, 86.7603238961461,
  13.5865545693098, 4.95627940006259, 61.1583587698066,
  13.9585752430574, 4.37130749064627, 61.8790587652959,
  14.1158877937273, 5.80332041778817, 61.1101109530874,
  3.71485169993295, 18.1102556966989, 59.6482905184618,
  3.02128279270173, 18.4612635983734, 60.2773816278285,
  3.91846415341326, 18.8029475757733, 58.9563946235094,
  15.5625795867826, 7.83360061471947, 82.3608626843385,
  15.3126473983664, 7.42832097083809, 81.4814979639586,
  16.1200949608325, 8.64912350193044, 82.2056240675801,
  3.82247061350724, 5.9422691325601, 69.2517075181748,
  3.50396472232506, 6.63686444994935, 69.8967589442977,
  3.91427295910467, 6.34867885032903, 68.3426401550791,
  28.0889432537582, 6.22627984084838, 72.1981165378426,
  27.4258704033709, 6.08863153032911, 72.9339068188945,
  28.2952904024379, 7.20108351688259, 72.1133896387968,
  11.5622919277592, 17.9446791005478, 83.54515201111,
  11.8972847672415, 18.6115561136894, 84.2107756636637,
  11.1674886535323, 18.4249271962654, 82.7618946196866,
  1.70880315699884, 2.72962190274191, 92.4392035748222,
  1.25038240668451, 2.23185856217449, 91.7029413440454,
  2.09222475970384, 3.57981818985675, 92.0784347458537,
  2.33226399398277, 28.1739401705963, 83.4204879379026,
  2.8320691918441, 27.5316500970239, 82.8394042730305,
  2.77231806502252, 28.2242425382635, 84.3170491942418,
  30.1307736973707, 27.2653644964995, 63.9147178431862,
  29.585244502228, 27.7333215158967, 64.6099977330463,
  29.6194351469867, 27.2328548761401, 63.055953608093,
  12.396000789532, 15.0959461772172, 75.8719381468277,
  12.887035955172, 15.5558407365722, 76.6117904701872,
  12.347518580698, 14.1155605474264, 76.0629708464539,
  21.2782906920176, 9.72732624908679, 91.6858108388381,
  21.5144409060003, 8.7914298851213, 91.9472129665113,
  22.0061309404257, 10.1078079859883, 91.1153003475395,
  18.1338787723882, 2.20582112233515, 63.5544476474892,
  17.3490385852415, 1.59888900712986, 63.4293105699623,
  18.9754798950788, 1.71172465859186, 63.3363278757986,
  29.9364417324311, 0.214126675930733, 72.4722356530209,
  30.5907653218126, 0.266987736770833, 71.7178707886311,
  30.3506827067146, -0.276141725139094, 73.2390741693574,
  25.5779936607684, 28.0170863612097, 70.1179938315458,
  24.6362311590477, 27.9201852475664, 70.440008682954,
  26.0019180264316, 28.807364781589, 70.5604281775001,
  -0.322391188502927, 27.0336040668785, 59.3791101384463,
  0.548741725526838, 27.5050516525526, 59.5164586734081,
  -0.198346832007921, 26.2881190887524, 58.7242321765252,
  14.0598293579625, 9.99599801481496, 72.8090485820983,
  14.4529897478881, 9.40435773813593, 73.5128857016116,
  14.5856637152384, 10.8448836294613, 72.7552764521902,
  9.72826869797064, 26.2178081011633, 81.7590742562049,
  9.55856451990728, 25.2464730125768, 81.5926151392165,
  9.06276380612131, 26.7643705271226, 81.2507704558511,
  22.1399709592699, 22.5768640067273, 62.0221237023795,
  21.8600329890327, 21.8260582722055, 61.4238549652483,
  22.2575899698015, 22.2342685953608, 62.9542149814247,
  10.5869429469486, 18.9592471860192, 71.887722380062,
  9.84126366487338, 19.625396264588, 71.9021381147237,
  10.2174800581782, 18.049352020338, 71.6990746626327,
  5.45373214354091, 22.689862840764, 91.465488461986,
  5.14840782391397, 21.7496362953578, 91.6163231501643,
  4.66890163600661, 23.3074614773416, 91.5166059593912,
  27.1091523855975, 18.3708346994098, 86.9610458462315,
  27.603030051787, 18.3417690870306, 86.0920003692763,
  27.7628512616627, 18.339688528933, 87.7171593929265,
  20.7840583621346, 16.7453308163193, 75.4840688923301,
  20.3920993316662, 16.4060243756727, 76.3391941800921,
  20.3828731693005, 17.6342719936545, 75.2630846750462,
  3.86203714151241, 23.2218110010577, 74.7976451122072,
  3.77698984697542, 23.2741390503674, 75.7926469880584,
  4.45175172489153, 23.9617876284421, 74.4741156683003,
  4.6492003943311, 14.4896904264417, 84.3309040144901,
  5.38775786845237, 14.6820483905562, 84.9770706114768,
  4.95116982398107, 14.7116814926891, 83.4037932174096,
  12.5504137786472, 9.89718069954809, 75.8201561566585,
  13.3116347772525, 9.27599274022483, 75.6339624122035,
  11.9248556013269, 9.9010746007381, 75.0399883514261,
  18.2274189878982, 6.88664913321818, 62.5911993349318,
  19.1911042112961, 7.0108228585292, 62.8276135395538,
  17.8569618333439, 6.1092762455187, 63.0995819566935,
  18.2711502844191, 8.25132921280715, 67.1160136945011,
  19.1849664234728, 8.46156675084586, 67.4634906600748,
  18.3141267961795, 7.43804949822536, 66.53573003517,
  12.982482096769, 11.0452102809762, 86.1115178331125,
  12.4638677906512, 11.7472449486776, 85.6234742624805,
  13.4018989663335, 10.4216055037076, 85.4518159524933,
  30.2373281760281, 14.2795042806639, 75.4095408678393,
  31.1162087658961, 14.7549648656031, 75.3707318363841,
  29.4962542604006, 14.9504133092313, 75.4358187475745,
  12.1329160737173, 3.60046175840295, 88.4830863776296,
  13.0379344176628, 3.3047928974759, 88.1772731637223,
  12.2166491823917, 4.4563632094213, 88.9934014495767,
  21.7846847098271, 6.61696161300294, 91.7037419959978,
  22.4684380006951, 6.95106414494866, 91.0550071230531,
  22.0472325420485, 5.70740005387556, 92.0258699301384,
  24.396240244761, 18.850638487258, 60.9464506937961,
  24.5134950646997, 18.1799588066846, 61.6788713879789,
  25.0006698266542, 18.6204479548051, 60.183773042818,
  11.9073997530759, 0.939963877668792, 61.4726285192635,
  11.7335914742636, 1.24866094924461, 62.4077738556775,
  12.7990970608273, 0.489280441591428, 61.4306719727615,
  20.952243763577, 9.83053769528038, 86.2964198657043,
  20.3706107369389, 10.1664191449472, 87.0372887300072,
  21.2223476677357, 8.88664684783292, 86.48645657022,
  12.329690027308, 6.14411790535259, 89.7077029066174,
  11.7308532342077, 6.93480825990769, 89.8349949269599,
  13.2701682106178, 6.39853628938575, 89.9330294975566,
  19.4005173858465, 17.7527402665406, 64.6998328518585,
  20.250509003462, 17.2286887139545, 64.7535377884612,
  19.5315762601999, 18.5396029718668, 64.0967817309575,
  3.45728280089315, 6.70256841259764, 66.2234032196128,
  4.40867851708954, 6.96606035304407, 66.0639723928479,
  3.00126964831216, 6.55314967384971, 65.3460628950043,
  9.84913147354695, 10.7612169643927, 79.9009934924933,
  9.79300112733357, 10.4343855374451, 80.8444078249015,
  10.1538784734124, 10.0161651126433, 79.3076748561117,
  27.1033367284877, 20.546981999884, 60.4969096967172,
  28.0634785058462, 20.3419235559941, 60.6868539042106,
  26.6357923551893, 19.7127162207979, 60.2046720043453,
  27.6548838969887, 11.8335878568926, 70.9752555086505,
  27.3931021240116, 12.0331279519032, 70.0309811556047,
  28.1323337518248, 12.6222757956899, 71.3625705888018,
  4.02083175278648, 28.1457881737432, 71.9410316125234,
  3.35602150661186, 28.6219834101842, 72.5165882416852,
  4.93490093027137, 28.5124698981536, 72.1143003395214,
  7.40313807884473, 1.83372138620403, 64.1225822172815,
  7.83176672831112, 1.71786041745418, 63.2265611702201,
  7.19712725184311, 0.936053005252626, 64.5121345462416,
  11.0039808934089, 9.62133397281773, 82.9368130901708,
  11.3524697236164, 8.68572789865953, 82.9933534228446,
  11.7598646645396, 10.2476420160964, 82.7460830205287,
  7.2573703988512, 31.0092131287819, 76.6309888111179,
  6.29980001977257, 30.9829466505149, 76.9179888829483,
  7.50827488237991, 30.1299113142104, 76.2261737187159,
  -0.103355749481144, 7.99963761701333, 71.4015966537979,
  0.8315510204592, 8.09628709041844, 71.0601172095992,
  -0.194677880411671, 7.12662050274646, 71.8806596836796,
  8.35941475276385, 15.4022201809511, 76.8309096041017,
  9.33085969372971, 15.6120544051175, 76.720165190968,
  7.81202560370813, 16.1568749457479, 76.4691620326303,
  7.94707428945413, 4.70293383831056, 90.734865944085,
  8.01139987700691, 3.7050586712234, 90.7452278790756,
  8.69966313020924, 5.09102595116386, 91.2668382635828,
  16.4585402488836, 4.07679207190117, 86.1180975626403,
  16.0026998996239, 4.81909764425683, 85.6269845275491,
  17.4476134068136, 4.15071229756241, 85.9905433055549,
  30.3454692447894, 2.8779604415952, 67.0853081645409,
  29.8179428873339, 3.57371316911395, 67.5727956867812,
  31.2282438080668, 3.25987132547798, 66.8117151324618,
  20.6718662462269, 10.6852153109886, 68.6797327901363,
  19.7258150942915, 10.956785717788, 68.856471954083,
  21.2500064486766, 11.4999992064686, 68.636361025383,
  8.27504887653133, 4.63505422798133, 64.2524226555542,
  8.28253294661343, 4.5683752535398, 65.2501690677565,
  7.72270317087211, 3.89285994073805, 63.8728678355042,
  6.99912466625028, 12.3301338970699, 79.0049416386455,
  7.11146477149994, 12.5364851237379, 78.0329339884672,
  7.66762448607901, 11.6384876336479, 79.2783158093043,
  30.9293758768568, 16.001189067435, 69.6833248841237,
  31.5658833516085, 15.3135861143071, 70.0326963389321,
  30.0305692224603, 15.584626856162, 69.5468605219193,
  2.92203334339994, 25.5848820133538, 67.6274285829131,
  2.21068300216736, 26.2845866385955, 67.5611403528595,
  3.82025614781735, 26.0238223556113, 67.6503887563306,
  27.620390563966, 26.3316078047216, 72.9680732132203,
  26.8852572876926, 25.8268178814967, 72.5155622194024,
  28.4583150923561, 26.2562656253283, 72.4275123556599,
  0.567750850246448, 23.7158535043579, 77.708366988372,
  0.174530455648181, 23.8526156932699, 76.7991509387139,
  0.169065464463156, 24.3745205417854, 78.3464952646373,
  24.6190010480547, 28.0694585012452, 75.3304461622765,
  24.1723552209798, 27.2354830726206, 75.6544716082018,
  25.6094760417064, 27.9790548658056, 75.4343040924017,
  18.7820754624663, 18.6292898623562, 67.8986735071234,
  18.7526252717873, 17.7559951870534, 68.3849749530978,
  18.344736686914, 18.5281439049724, 67.0050828342181,
  12.3233007445071, 21.2082152189065, 75.4948372293278,
  12.4097219290971, 20.2916158401707, 75.1044823167735,
  12.3733762023731, 21.8881598623399, 74.7632856382655,
  14.6176303730822, 21.5007600684469, 72.3303822377802,
  13.9022750723885, 20.8700346777883, 72.6311350853944,
  14.9852338193278, 21.9895894870828, 73.1215291936516,
  7.62173044260456, 1.17697592223645, 73.3167296441356,
  8.24832465876366, 0.772727651340962, 73.9830351474552,
  6.77837808577791, 1.45365064144384, 73.7773899332712,
  -0.129383504648538, 14.6042524459504, 65.447455158437,
  -0.451137464133561, 15.5496708380632, 65.4990153505488,
  0.859600151829637, 14.5963047298062, 65.2996439239954,
  24.1207448958887, 29.5649554933352, 68.2494224351414,
  23.2951957833838, 29.1761533015686, 67.8403973521455,
  24.5511839412022, 28.8844862184378, 68.8424517718443,
  8.13369075861067, 27.5882910362941, 71.7169622515939,
  8.077483354452, 26.8413845549812, 71.0544130565218,
  8.87271834206864, 27.4041462392633, 72.3649814832643,
  3.26256556433436, 6.47256284534099, 89.1882323413804,
  3.84955147020241, 7.23114823253915, 88.9053971302739,
  2.89976803603863, 6.01185246999264, 88.3782175862624,
  21.1366468490824, 13.7491463017756, 54.8812006409547,
  21.009335524458, 12.996672821669, 55.5274014521262,
  20.6810772072928, 13.528583291515, 54.0187574486316,
  14.6348563370127, 25.1641627228708, 89.1115007453077,
  14.6171643345712, 24.2099444807812, 88.8129131710301,
  15.4445964015767, 25.3216060911051, 89.6767729042178,
  9.70289952891882, 7.13936502529509, 56.5639736999227,
  10.0248110741827, 7.92155993848978, 56.0305469713103,
  8.8267892341267, 6.82467917111945, 56.1987291728713,
  24.7802211001246, 3.74235492934249, 84.4259036786186,
  24.9171183348934, 3.37953837463356, 83.5041535526398,
  25.6284324069498, 4.16279938903955, 84.7480279330361,
  4.83413509423501, 13.9337538542197, 74.6340143542237,
  4.83889500026979, 14.0691402615443, 73.6432329131348,
  4.55391302262368, 14.7811998925328, 75.0849143461613,
  29.8486045425795, 20.5259341396683, 61.0200595275854,
  29.9812054592859, 21.2779959505323, 61.6656755353861,
  30.2084656067541, 20.7879589838245, 60.1246026634451,
  22.5056262253389, 26.1013962297476, 84.2079096807423,
  23.2792666650721, 26.4935943667078, 83.7102540856021,
  21.9797271693794, 25.5114243139883, 83.5952406660564,
  16.9618347073679, 18.0125204615046, 80.9495697217588,
  17.6849755497321, 17.4232047442446, 81.3098117341548,
  17.2943128135903, 18.4884105460697, 80.1353296243088,
  24.3885539319905, 23.9555350088271, 66.4102234135616,
  24.9797352895296, 24.5483527281191, 66.9570979459654,
  23.5905932845344, 24.4734130248373, 66.101903505601,
  26.3954421911863, 14.9488560225518, 71.8897147664199,
  27.2307422477328, 14.4031134775988, 71.8230897698963,
  25.8625739020554, 14.8466183255054, 71.0497154570504,
  12.4498108121183, 25.2590427505211, 72.0773386874335,
  12.6368463489401, 26.2253838169532, 71.9006959652718,
  12.786135617029, 24.7092290107715, 71.3127535207029,
  1.08076495034946, 25.7884603475024, 74.8570327415817,
  1.42549232498133, 25.654367826259, 73.9279567312758,
  0.413315787844941, 25.0752404759122, 75.0711099011314,
  4.35854600977722, 17.306671095722, 70.8481166714017,
  3.72090885167802, 17.2637140809047, 70.0789784851899,
  4.83660333820836, 18.1849181107947, 70.8361428980094,
  4.01461558985599, 30.9272555011578, 93.5845612581623,
  3.04675916307518, 30.9764013117621, 93.831216131293,
  4.45729094498604, 30.203767467981, 94.1142815577643,
  0.753173735665025, 8.43823819772177, 89.6863621995417,
  0.0524844150499072, 8.42151432620373, 90.3996326868727,
  1.38439989007266, 7.6744499687357, 89.8211994468218,
  18.215903105152, 27.7687438324957, 82.8840733166946,
  18.3008258881755, 26.9054675390899, 82.3865372253735,
  17.3821279160995, 27.7547672058028, 83.4360004749563,
  6.99087073384816, 13.0545922636037, 76.146251420922,
  6.09339081928903, 13.1371553422208, 75.7129926748912,
  7.36228164677989, 13.966643692963, 76.3200792781798,
  19.2714891467567, 13.6819756851126, 59.433654977521,
  19.6963411780748, 14.5813528635834, 59.3305945955555,
  18.9149096343011, 13.5862741721088, 60.3630054344024,
  20.6822453168831, 23.3611778950067, 78.4570982526248,
  21.2709655736981, 23.9109172340822, 79.0497154294672,
  20.4998627506587, 23.8621439185549, 77.6110665494436,
  26.9331001113161, 30.0158901157124, 71.076601230855,
  27.0000821191062, 29.938015180025, 72.0713116937658,
  27.8393879955545, 30.1968129439839, 70.6946206016433,
  17.2767203656058, 25.7784967356587, 90.1122556081651,
  17.8318952963873, 25.5954113734387, 90.9235881826206,
  17.7334512623954, 26.4622589296401, 89.543163216721,
  30.5975081991643, 23.9959719114518, 83.0604116858222,
  31.4930190664989, 23.871462779771, 82.6331438978794,
  30.3991768732375, 24.9728510216862, 83.1402357996208,
  18.7594794621472, 2.69982581398044, 89.6527453416839,
  18.2459688769234, 1.9161511404894, 89.3032301274344,
  18.5938971304764, 2.7959412456556, 90.634246393763,
  27.374426076891, 23.5632767373968, 75.46687971609,
  27.2080562769593, 23.4876529053242, 74.4837204585465,
  26.5469225335118, 23.3057100337101, 75.9657757762537,
  4.45025654692929, 0.659081663576113, 77.714831579859,
  5.05299172532584, 0.624750091151799, 78.5120339681257,
  3.66196629115152, 0.0628938299103424, 77.8670108807995,
  15.2717286661362, 4.70514011142396, 75.4257789465738,
  16.2445268441042, 4.89803568852626, 75.5540559954816,
  14.9576181082917, 5.12679649375496, 74.5751671357634,
  14.6858710573616, 17.0746664465142, 59.1129262562239,
  15.1884077959833, 17.9391237792602, 59.1259779303391,
  15.3324886004809, 16.3140241911952, 59.0554013715778,
  23.9075707300587, 13.9216337107003, 59.5566636178039,
  23.6774289529867, 12.9561434344179, 59.434748529114,
  23.1426717014669, 14.3939065231696, 59.9947136910394,
  20.856458810072, 29.4380128521897, 80.2727852499043,
  20.9185095175549, 29.7903387948028, 81.2066032942056,
  20.8431535972118, 28.4383238820004, 80.2938787131687,
  10.5847284646343, 2.57992120708627, 69.5979816734372,
  9.61410052929525, 2.4744408000038, 69.8142114004894,
  11.068455713284, 2.9317420962041, 70.3993742182579,
  10.1566909391021, 27.4366649886751, 74.0036436842253,
  10.8552304171317, 27.548361734588, 73.296843546572,
  10.5238279158964, 27.7338074685432, 74.8850725168193,
  16.4888934535359, 10.8323737854984, 76.0438493104859,
  15.9262501535924, 10.7424853850133, 76.865647699683,
  16.3321326444525, 11.7286246724537, 75.6289271534885,
  21.4554078165888, 15.5424422105626, 63.800127271673,
  22.0831460354238, 16.1173896834511, 64.3248940122663,
  20.9452689729593, 14.9502911699802, 64.4239185070695,
  7.7464518179719, 2.42072064094099, 88.2963856740883,
  8.50370065347325, 3.0542416887946, 88.1375609812402,
  7.80779234662407, 2.05394520724072, 89.2246707169381,
  6.98993691526104, 8.31556756568762, 63.1276733310745,
  7.53312986812937, 8.79250427778859, 63.8186673893735,
  6.44923268785109, 7.59752638761177, 63.5659150509603,
  27.5179013804297, 13.4447139516522, 81.8333213649339,
  27.4121394910251, 13.6521847173585, 82.8058285906791,
  27.2862589406676, 12.4857297152369, 81.6699475163288,
  29.6033697143735, 19.69967329105, 75.4400075812739,
  30.1441832631518, 19.2605822803402, 74.7225678348341,
  30.1908765287454, 20.3050364015874, 75.9770096738835,
  0.234398319091294, 21.4920436677936, 58.6904938437271,
  0.63526902932804, 22.3736489422646, 58.4413456675365,
  0.877210325346038, 20.7588990172017, 58.4684766238471,
  8.39369799183905, 25.742434867288, 63.2737867054948,
  8.70923291963911, 26.6011513040755, 63.6775735187134,
  9.12838618429806, 25.065240013887, 63.3142884386492,
  27.4692800580396, 19.7613988337837, 77.0844288736663,
  27.576024703598, 18.9929514064499, 77.715375885759,
  28.2609475840632, 19.8047926837221, 76.4750197319336,
  16.6970390352453, 14.5797775079133, 81.4017266854373,
  17.6675224480377, 14.7505044846294, 81.5720623684757,
  16.1557027047488, 15.3343039807914, 81.7727317784089,
  4.87135786556505, 15.6881181224951, 59.0150414111261,
  5.86732462891872, 15.7356331125384, 59.0911500966752,
  4.48010587879956, 16.5913739710433, 59.1912536550696,
  25.0393206053834, 20.9863865841899, 62.6436280820761,
  25.9298460062997, 21.2938493760957, 62.3083205487335,
  24.6946773683361, 20.2565564404218, 62.0532307578908,
  25.7731027178197, 23.8430902250405, 91.2614558849752,
  25.727257242173, 24.6157614378941, 90.6283070958347,
  26.6144057513381, 23.9019126071441, 91.7988097098954,
  14.7518207917018, 3.4046887103926, 66.7726585101619,
  14.6961473930002, 4.35774621720276, 67.0702855609987,
  13.8388755130982, 2.99688548899399, 66.7877399852973,
  24.361341713538, 20.645890483452, 79.0089159704995,
  23.5822362842993, 20.6452270683806, 79.635808537062,
  25.1907895667902, 20.3945347356405, 79.5077511604947,
  1.34613989321356, 18.9177822132864, 61.2216049859388,
  0.711702448376721, 18.4510971738072, 60.605411670075,
  0.932778477987554, 19.769779622829, 61.5429035301854,
  5.61014603648751, 26.3492458101822, 67.6551852659054,
  5.64433169095194, 27.3471878447386, 67.7094350280623,
  6.10391205055807, 26.0425339334902, 66.8414758902405,
  -0.0717086968810548, 20.990781275429, 77.4351476910271,
  0.754783077131679, 20.4399924234082, 77.5515220351882,
  0.147530212612323, 21.955615268636, 77.5801637801912,
  18.6632756199927, 22.3381662915204, 69.3865597512632,
  19.0690946846627, 23.1350546723533, 68.9390334445012,
  19.3117930116174, 21.9608774758069, 70.0476787589296,
  17.4228684139651, 28.806232661545, 79.6439388206473,
  18.2132812999347, 29.3356721058475, 79.9520643543342,
  16.584766363921, 29.2229699837278, 79.9959543856607,
  26.6631336076014, 3.94977905418937, 87.9122939413125,
  26.5813978463765, 4.79960576280398, 88.4329798645544,
  26.8109699993122, 4.16340708625219, 86.9466296801933,
  9.80632137349007, 21.003978145478, 76.8456702677399,
  10.7814100925068, 21.0938633600236, 76.6428830929671,
  9.31026900904261, 20.7825274930268, 76.0060920044106,
  28.0333291801266, 28.0186675743656, 77.8178353018907,
  27.8945359632961, 28.9669375222964, 78.1033533377714,
  27.5112026775565, 27.8419368994342, 76.9834791526043,
  10.7625872319892, 15.2941216222828, 85.0287442460609,
  11.2731977776605, 15.6713807238674, 85.8013712200404,
  10.8127386416145, 15.9262468140779, 84.2555026421553,
  12.1334344708687, 16.203797497322, 87.5476671757727,
  12.934381822502, 16.7048149134197, 87.219848798194,
  12.3796616439432, 15.2473279090089, 87.7043136116462,
  5.53877518683474, 23.0035254489704, 79.7579261956955,
  5.68659201692072, 23.0899196612364, 78.772692099234,
  5.85090997937729, 23.8357929396173, 80.2160775847546,
  24.9371983314782, 9.32459139382173, 60.7826885169432,
  24.5941074757849, 9.02818210762627, 61.6739966565878,
  25.9154845235257, 9.52047479661333, 60.8504071920644,
  5.57639999752779, 15.6160352094201, 82.0398544098395,
  6.29772476247566, 15.1773629866646, 81.5038905449609,
  5.96269891673037, 16.3804235283633, 82.556074946903,
  9.06361450565748, 20.1587908142875, 67.8699584926229,
  9.55102604390856, 19.3860470548093, 68.2765259219225,
  9.51701401735302, 20.4293283762049, 67.0207009872772,
  19.9662647021786, 19.901487592459, 75.2470357011047,
  20.8714483285809, 19.9889007265041, 74.8311011551847,
  20.0458193745383, 19.9890770985217, 76.2400105912874,
  14.7665393285821, 30.6289815614142, 67.8006096673321,
  15.5126827069501, 31.2385670797344, 67.5328867606322,
  14.377797682335, 30.9390171933749, 68.668225849401,
  17.5272077287286, 21.9265856424685, 66.9558878277129,
  17.9139914124103, 21.8325174378504, 67.8732479287188,
  17.4051183053097, 21.0203774931416, 66.5510656904937,
  28.3361109086436, 29.3143632211966, 64.7416286534783,
  28.3803276153796, 29.8578144064833, 65.5799040808027,
  28.0470211004929, 29.8966126247407, 63.9817518773521,
  0.844698326477473, 28.4820643050413, 70.2366753074504,
  0.925464732386518, 27.9532725242496, 69.3917752895526,
  1.68221960995381, 29.0089167123226, 70.3815360704819,
  29.2281980220963, 3.83564524817082, 91.3665524453048,
  30.1823661325185, 3.80414704268867, 91.0689435070908,
  28.8307629557167, 2.91980042840347, 91.309336764612,
  6.27597771078518, 0.918949036443961, 79.8207831293276,
  5.67183075148217, 0.387000664927161, 80.4141105108005,
  7.22821352907001, 0.740538077612613, 80.0686066071183,
  9.37652853214227, 16.3666675388686, 79.5421048842055,
  9.53911124202632, 15.4528440210703, 79.1699578154739,
  9.95241124032949, 17.0290471529699, 79.0629260519998,
  26.4443454903036, 7.01145990771357, 83.0435018585051,
  25.4643686703635, 6.854381693852, 82.9211422773109,
  26.6426894005501, 7.13920837355426, 84.0152734483056,
  28.6056554349836, 10.6285033151973, 64.1478832063673,
  28.9601118600496, 10.6462320029135, 63.212978753302,
  29.1300511252003, 9.97258262290964, 64.6908170932365,
  5.26284949259946, 19.9579677202708, 92.0226545156126,
  5.92080008040872, 19.3877692072874, 91.530745296556,
  4.6863587421917, 19.3795069036229, 92.599751992905,
  19.0332381384945, 16.3057945707548, 69.456672738175,
  19.1517555549889, 16.0868344543881, 70.4251819479547,
  19.8053662429288, 15.9418769182222, 68.9357292359428,
  21.7618438731172, 18.8474633575518, 84.4368054286931,
  21.7094447552729, 18.3641217619463, 83.5629431773018,
  22.4041526987989, 19.6098540330216, 84.3580664268698,
  25.2064403681292, 8.20222270771618, 63.4723447480283,
  25.6745115321751, 8.73971673934853, 64.1737786731761,
  25.065420021642, 7.26998193803255, 63.8055720116432,
  16.3144614193196, 2.09015911433849, 78.6937899233089,
  16.6815954923491, 3.0185427019518, 78.6362009775724,
  16.699399479541, 1.53322146387351, 77.9578258322776,
  16.8983583499059, 29.1169192300368, 66.5951228685976,
  17.5100404041583, 28.4609564800243, 67.037342197779,
  16.3628803153503, 29.5950776660542, 67.2912749960624,
  24.013548931869, 8.79542964498769, 78.4466658478851,
  24.072859852344, 9.66703153204646, 77.9600526902455,
  23.9792685728413, 8.96517449396963, 79.431557488234,
  1.46843506946256, 11.5893020834602, 57.4343039891899,
  2.19825175298284, 12.2662280553643, 57.5299012538845,
  0.705247095400254, 11.991144994141, 56.9282739590709,
  14.1244731952609, 21.7263952648853, 58.2278692835717,
  15.0010677960121, 22.1346267096248, 58.482680965917,
  13.3817891490068, 22.2269554107667, 58.6726837929966,
  0.272245107796799, 20.5339589409414, 84.2269263555174,
  0.0814549861655429, 20.3179975299226, 83.269346176922,
  -0.077964063553619, 21.446293425273, 84.4390567988803,
  7.77266753813813, 8.14950606982496, 85.511509421343,
  7.52786491373968, 9.11838899232532, 85.4749367871091,
  7.00238510464333, 7.62449620261803, 85.8734895478481,
  3.61218707225448, 4.97308336842853, 58.5798111850477,
  3.52793440424236, 5.44703212913148, 57.7032987435154,
  4.52996730207121, 4.58455400141445, 58.6618135065099,
  2.74115456498723, 10.1595850335472, 80.5348487326313,
  3.16866552153609, 10.4855794537918, 81.3780343705546,
  2.7285576122979, 9.15966716781351, 80.5324868330868,
  3.08843467346227, 27.8729247981015, 92.6745668560774,
  3.53350569664363, 27.5285641296458, 91.8479305912396,
  2.24917641582167, 28.3558787731994, 92.4247648646537,
  1.02291762213251, 12.050775627545, 61.8642221205671,
  1.28110991794552, 11.2546674426074, 61.3169118828973,
  0.0274993556241873, 12.0853833603856, 61.9533556133137,
  19.1804075961343, 25.0274194727632, 82.1555497876227,
  18.8174191904336, 24.5499526989333, 81.3553842439911,
  18.854309261663, 24.5789020388067, 82.9877108223343,
  6.50631317589722, 8.29692669291425, 80.0516549105519,
  5.82197133320795, 7.63177651267426, 79.7529050485079,
  7.28189787800878, 8.28357809521215, 79.4205525537271,
  12.5061311873758, 11.3666437876874, 65.9064613637445,
  12.0177321320997, 10.4982981080923, 65.8201935045268,
  13.2102284557224, 11.4248202047576, 65.1987449366329,
  2.79327416250389, 22.9654994136934, 82.6172819138536,
  2.95060327963143, 23.7130031961618, 81.9719249241965,
  3.66529361257169, 22.6780697269675, 83.0134715829416,
  1.66851457205825, 17.0393776028227, 75.2405245129476,
  1.08980742557374, 17.6191164687714, 74.6669385246981,
  1.37455251631416, 17.1137533719943, 76.1934434784126,
  3.02634580459589, 29.3350770896225, 87.1410525948064,
  3.54026559661165, 29.6926175172987, 87.920829030685,
  3.07310513002204, 29.9867121930473, 86.3839626018266,
  14.1936373174412, 19.1567579869002, 81.8529335140877,
  13.5081669564744, 19.2086786035091, 81.1266865631082,
  15.0588282613145, 18.8306644541318, 81.4720035487054,
  8.79733670818162, 15.2338159719895, 62.3303966333837,
  8.80460963452538, 14.2338677934353, 62.3375201682096,
  9.22323832347504, 15.5642752686787, 61.4881351138293,
  1.23630445265045, 23.9505571665065, 87.6202172573987,
  1.50868869060006, 24.8964365427496, 87.7966231317751,
  2.03290836831381, 23.3524225006904, 87.7077222463932,
  25.8611803845043, 12.3406943482734, 54.3005875818978,
  26.698882805436, 11.8425534945353, 54.5244409799114,
  25.8688562525674, 12.5872935583249, 53.3315004286182,
  16.8286643009966, 9.48691321055162, 63.6287351063199,
  17.023873095435, 8.53437047233287, 63.3951631507246,
  16.5293672155599, 9.9763692307903, 62.8096782957742,
  18.073919582173, 18.193113538273, 59.8649424061281,
  17.3023271460463, 18.8239810430805, 59.9464979325509,
  18.037924777474, 17.5246623181573, 60.6078268792196,
  4.39278631499144, 27.0328924500298, 90.4493528999234,
  5.01967871992643, 26.5114991931655, 91.0282786156515,
  4.91703670952806, 27.5594827144737, 89.7801263185467,
  16.4068180102142, 28.9592408410082, 91.3646342630332,
  16.2516770598453, 28.0536243755822, 90.9699317129174,
  15.5271434963458, 29.3953171423753, 91.5543978239092,
  24.1126509462335, 11.3684084891278, 74.2198570056158,
  24.1724647458329, 11.4676499975219, 73.2265929760702,
  25.0162831312509, 11.5101335576227, 74.6240387458773,
  23.8842974596039, 9.51832537895201, 81.3040526685208,
  23.1149401949332, 10.1056512735812, 81.5553248173882,
  24.7307152053288, 9.90114423391991, 81.6742238775622,
  15.602536828458, 8.49878973566253, 78.6095811941131,
  15.0324601233133, 7.68856341597843, 78.4733980044657,
  16.424135422988, 8.4271912174814, 78.0440288962126,
  30.2161133500984, 27.5498111266558, 76.0256610294657,
  30.9990331870341, 26.9392840805964, 75.9061066277795,
  29.5951491934154, 27.1657018679835, 76.7089352010228,
  30.2983283936525, 10.515728666126, 67.627134323001,
  30.2590950925116, 9.83578993159223, 66.8949157317578,
  29.6003206611863, 11.2145575105092, 67.4708542805279,
  6.51790638196642, 18.8914951471406, 67.7019297766848,
  7.28892222783487, 19.4893189264528, 67.482518531967,
  6.08046963740129, 19.207106754848, 68.543973960552,
  19.937013262135, 10.4001203553615, 80.1076883691582,
  18.9712041909555, 10.5736943482064, 80.3002627886307,
  20.1576953133171, 10.7270767990162, 79.1887765582434,
  28.8677358242841, 10.7713709646829, 82.3766128880841,
  29.719361753627, 11.2869623777033, 82.2822795891356,
  28.8260815648444, 10.3602550484045, 83.2872437826035,
  19.1220513292712, 10.9685031486476, 88.235390551092,
  18.5110169724673, 11.7600418817657, 88.2455615283796,
  19.0007328768911, 10.4428958486425, 89.0774230916113,
  7.84937531752638, 12.5868925895794, 65.1599772478751,
  8.51046430399651, 13.2163031246313, 64.7515611238867,
  6.92619981100869, 12.9548984640569, 65.0489877865921,
  23.3431155228062, 20.9919074338768, 84.7704919367026,
  23.0643219339707, 21.8955594782596, 85.0955874880518,
  24.2972989184597, 20.8274697354142, 85.0204805180089,
  28.7038893262137, 7.99379727553314, 81.4987376820394,
  27.9946496222388, 7.58295919733997, 82.0716173516143,
  29.054047777027, 8.81891600148483, 81.9420977472323,
  30.2998333791162, 23.8209183859305, 75.1927793479139,
  30.4373277350678, 23.5372046400677, 74.2437789198371,
  29.3892017367158, 23.5402154734852, 75.4960216385066,
  27.4734256892574, 11.1128818688144, 60.5364811037804,
  27.136785972167, 11.4268047740321, 59.6487164331289,
  27.7649656198748, 10.1590628528228, 60.4641364178081,
  16.2815404922872, 13.2773258262232, 68.4800475320445,
  16.6786726545759, 13.8750767149553, 69.1764525296543,
  15.3665554146488, 13.6037959213605, 68.2429408373266,
  3.90983378790478, 12.6760724299582, 62.2541155044809,
  2.95177932220319, 12.561205678144, 61.9915564252685,
  4.49682737641748, 12.4744631891615, 61.4700286208575,
  5.1695861862238, 9.26153957398261, 86.2216290094014,
  5.89247340044758, 9.89949710109703, 85.9562156165407,
  5.1564711444019, 9.16806076091416, 87.2171638943679,
  8.87360644521947, 14.6256619677677, 73.1229692710886,
  9.40656944405837, 13.910589105587, 73.5753200681934,
  7.91285214971698, 14.3510287030346, 73.0838827826872,
  27.2849333388371, 9.14918874154237, 74.9419725882668,
  27.7597079523974, 8.97864280485422, 74.0785473455284,
  27.5084537329657, 10.0671636514025, 75.2696320124802,
  28.3933078070397, 5.90350139955838, 59.1453186657329,
  27.6652885100541, 5.6287078013777, 59.7733922136678,
  29.2529199163593, 5.47489080769985, 59.423455290538,
  22.3545334251534, 12.7634939755702, 68.7380791373609,
  22.4546221877372, 12.683196861841, 69.7298122734067,
  23.2583291109152, 12.8392756323748, 68.3168778803706,
  16.0705901145794, 0.297539015945581, 76.1856792408459,
  16.9027650803026, -0.158394051239547, 75.8700689357689,
  15.7758686319277, 0.96446788727604, 75.5013217843589,
  19.6064449647197, 29.7789873259829, 73.2980960604531,
  19.42532812109, 29.001321549799, 72.6960722822633,
  20.5656536629979, 29.7656322331758, 73.5804793365933,
  7.29050523279844, 11.1131945230557, 85.6625780624524,
  6.99712696616695, 11.7370138843086, 84.9381620237051,
  8.25511372544991, 11.2746124963252, 85.8710839228262,
  18.4199429507174, 27.3018679448616, 88.0717215845263,
  17.4618630852654, 27.1770082366264, 87.8138591702917,
  18.9615885355978, 27.5017043748249, 87.2552134941566,
  25.4980089800706, 1.68054408969872, 71.5657349067315,
  26.0507979799142, 0.894239924019981, 71.2897818660014,
  25.2414641240284, 2.20829936717413, 70.7560071105338,
  1.46773213462562, 15.5979889453204, 59.2581899047403,
  1.83205596942814, 16.222518041993, 59.9490093824652,
  2.16592057766443, 14.9240189819434, 59.0167413875102,
  21.8040729656955, 7.18458682528768, 78.0524594025881,
  22.6464519940204, 7.71925993063639, 78.1197070274917,
  21.9974080862394, 6.3132562937599, 77.601455371573,
  8.20783766029385, 9.51913613568503, 71.7201326491344,
  8.76857404327345, 9.92671463219946, 70.9994007447608,
  7.82399479713381, 8.65479074063702, 71.3952146680062,
  12.6918566748482, 5.34072507074518, 82.8335542203949,
  12.5717884752071, 4.35849115885115, 82.9777768599501,
  13.4040738427615, 5.49240289368814, 82.1481780143906,
  1.57972515850074, 30.3866351789937, 89.4921827833009,
  0.611566344491138, 30.5302251171307, 89.2871207426368,
  2.11626313840173, 30.4859875722146, 88.6541755649042,
  2.10505184736816, 4.95365249774944, 77.5720148655197,
  2.26325730078292, 4.12803175297301, 78.1136064277737,
  2.92359960038345, 5.16346696983466, 77.0372649582386,
  16.7617653371212, 16.6984118872123, 65.2082200695842,
  17.7198929776989, 16.8951199815888, 65.0001399168356,
  16.2392089648999, 16.648707790645, 64.3570653594196,
  30.043848603907, 16.6460027386616, 81.6388425268079,
  29.8496718163208, 16.9566689830003, 82.569316524183,
  30.8442156297418, 16.0465587080695, 81.6477575783464,
  11.5932066801101, 8.85815382385389, 78.2722703428694,
  11.7567924141382, 7.89352776036452, 78.4789978573891,
  11.8690665488205, 9.04859481565048, 77.3301272743928,
  1.38651374387345, 22.2678197397492, 73.2825224892886,
  1.1613750931835, 21.3206402421111, 73.0541289972194,
  2.0010409981592, 22.2834953510866, 74.071262325324,
  16.8899059711919, 0.649990055187679, 89.5971620172808,
  17.0755774184927, -0.0722143407715627, 90.2634554392161,
  16.864010124551, 0.256913874210877, 88.6780208305878,
  28.3098356594146, 1.76710219968168, 68.9219561831521,
  28.3179123737593, 2.72359467018124, 69.2136013795175,
  27.3646565657844, 1.44875099289745, 68.8492307398501,
  8.09814217512077, 17.8017473473274, 61.782423247866,
  8.98896877715635, 18.2560163387738, 61.7741983760739,
  8.17571285283402, 16.9244000328509, 62.2559678389447,
  27.5397319225729, 6.01702947777752, 78.3046823129167,
  27.2310047760707, 6.34470573323956, 77.4117568845528,
  28.4962378650769, 6.27451842707209, 78.4417801719287,
  29.8092697222482, 27.9842915977131, 67.2360738632227,
  30.0441700846757, 28.9512538779248, 67.1370497834279,
  28.8383521845128, 27.8547971881517, 67.0347027312046,
  7.88275814502351, 4.16841985996872, 84.9114107017594,
  7.40881325712087, 4.54441571786976, 84.1151674235635,
  8.73199290400749, 4.67409973189448, 85.063358690435,
  13.9418327629897, 29.8633840797309, 77.0072624505856,
  14.8913129110342, 30.1770994867812, 77.0156345380564,
  13.3354201925645, 30.6305848991622, 77.2162282303062,
  26.0767591433726, 14.802900694937, 61.1365093258999,
  25.3079927941299, 14.4186784226385, 60.6252642322885,
  26.0987429222519, 15.7946406390523, 61.0101424128555,
  7.81646381866283, 3.84832008003883, 67.0821959911745,
  6.84549149207687, 3.61342946301336, 67.1273528183178,
  8.21012561014931, 3.81679918904083, 68.0009107604878,
  6.25014388904857, 5.41517527167863, 82.9123233648633,
  5.47231145019796, 5.94916994408485, 83.2437240089687,
  7.01153807916791, 6.0291529481621, 82.7042120964695,
  8.69951162621349, 25.3294810556054, 60.4517882729975,
  8.59045513013801, 25.313942437601, 61.4457023698963,
  8.89437009814596, 26.2634982873024, 60.1523855562275,
  4.63635200385804, 25.955989259908, 70.1625204971076,
  5.22279920805934, 26.2617549115937, 69.4124624707298,
  4.01950161956502, 26.6973497344975, 70.4268692253324,
  20.4687304231677, 25.2947891988138, 68.2615363492777,
  19.5352145654396, 25.2871237804757, 67.9030821894025,
  21.1164139665391, 25.3681496173374, 67.5031668637102,
  20.4925851876261, 2.59240286838235, 69.9347225631718,
  19.5469658414012, 2.59509876940357, 69.6094583872119,
  20.6605186815551, 1.76102751123041, 70.464452076355,
  7.06554922555855, 12.6448767683767, 70.1045659636218,
  7.1538353436727, 12.0348660668346, 70.8920254897896,
  6.11558065947085, 12.6507109589245, 69.7922749364277,
  16.2423616187034, 29.5130687480783, 70.6829534306786,
  16.944695124421, 29.8442079334449, 71.3130918969392,
  15.4590439007081, 30.134443161061, 70.7004803118944,
  10.2581665372297, 16.4630693410438, 74.9126362312114,
  9.70598082408289, 15.8432374985769, 74.3550526722172,
  11.071574079992, 15.9820242908205, 75.2396894822779,
  8.6429784044077, 25.1873769611663, 70.7304704166312,
  8.1938490732616, 24.3286046765249, 70.9770327962352,
  9.28886070888029, 25.0236597091378, 69.9847944077926,
  5.16047529609204, 1.5501297567117, 62.1651350809984,
  5.06178651655697, 1.97222465477008, 63.0662990071667,
  6.0075074335381, 1.01935454029644, 62.1366004043241,
  30.0091844428152, 16.8944148701636, 88.839916437383,
  30.7171139131802, 16.8708977420717, 88.1340249374519,
  29.7185115134871, 17.8395279829248, 88.9891493166109,
  14.1835830514531, 11.8523633264093, 59.1199232528496,
  15.0615385382979, 11.8166849369948, 58.6425123023594,
  13.5829190999451, 12.5094279765521, 58.6644357525914,
  12.4680213862993, 20.3616344857315, 56.3672410804441,
  12.9649374241859, 20.887063841441, 57.0578918195662,
  13.084712820771, 20.1348640919252, 55.6134063086657,
  22.9012772552575, 8.15487477162337, 89.2969723162933,
  22.2075233948852, 7.80225956766804, 88.6689849763269,
  22.8793825669761, 9.15461486956046, 89.290619427046,
  28.8179961003559, 14.517563547047, 87.269047165288,
  28.4758870871545, 14.1801686205107, 88.1460455043024,
  29.3725733707297, 15.3358707903572, 87.4201011514349,
  29.8683288031957, 25.3269650048596, 68.2370613354395,
  29.2102972343912, 25.0120883111257, 67.5530678250902,
  30.0425786490364, 26.3030944080486, 68.107414201054,
  20.1908002190034, 11.2194573719176, 73.4340060163058,
  20.9473328728296, 10.9290892424098, 72.848049795193,
  19.3243746683708, 10.9276249843869, 73.028863297256,
  7.21204532828502, 17.9364643933118, 83.0907470972552,
  8.00812616744361, 18.0153718001828, 82.4907229988513,
  7.43134469997089, 18.3202977711658, 83.9877307780562,
  28.204720728736, 6.25334474639828, 90.7608672119762,
  28.761743195374, 5.45120961546742, 90.9760536506452,
  28.3605269339906, 6.52211921820587, 89.8103490850009,
  12.0475148451367, 25.09302494948, 60.088319548379,
  11.2999787033775, 25.7142608183396, 59.8532542127678,
  11.8469806024476, 24.1803724612276, 59.7321574319264,
  14.7961035774128, 27.6707303006478, 68.4977486746079,
  15.2464849897548, 27.0666765884302, 67.8402719098679,
  14.8835437551838, 28.6192163186716, 68.1932351462964,
  15.1090396184581, 2.72385618705162, 88.0077248521868,
  15.6841891469903, 2.18274828247736, 88.6212436012372,
  15.687093201087, 3.3060581830215, 87.43597762526,
  4.81473241966652, 18.4585428716533, 65.6274042680737,
  5.25233296809315, 18.6459723683664, 66.5068222254629,
  4.75142188204685, 19.3054005393221, 65.099366517021,
  21.713270766104, 16.5977426284185, 72.7937335958786,
  21.3961370294633, 16.3984372727257, 73.7209356063793,
  22.0069920178732, 15.7498235494615, 72.3524161797258,
  12.3523120839158, 1.91683246425007, 67.5455065901048,
  11.861255579286, 1.8234055246042, 66.6794032959135,
  11.6973900120607, 2.07327852685183, 68.2848317616589,
  7.58671510327947, 22.4399527164155, 65.0551471641907,
  8.42220351650707, 22.8256999506892, 65.4465014571435,
  6.95093930572211, 22.2064294624582, 65.7908482074831,
  5.83932948814543, 0.752829429748427, 57.7289022658732,
  5.95608286896397, 0.266552697647748, 58.5948720043081,
  5.24126091717177, 0.22334454316854, 57.1272713663202,
  22.7964382983735, 24.8728197650631, 79.8006148750571,
  22.1254683952521, 25.5786700487589, 80.0277156590976,
  22.8819015434241, 24.2354183736945, 80.5663925843349,
  14.3007744817428, 11.6520119536405, 63.8202032350196,
  14.7064730300922, 12.4799522159427, 63.4330035321193,
  14.3229899375342, 10.9200395395885, 63.139231239567,
  9.37560604882149, 9.88094651277723, 60.8991798472524,
  10.2501731826952, 9.4395338336125, 61.0998965008227,
  8.63725491912658, 9.21191682567411, 60.9842497423561,
  27.8799831768594, 22.8901726001433, 72.7988022046362,
  28.7685325458238, 23.0546035682908, 72.3705003535695,
  27.6423180368084, 21.9226583236634, 72.7125966015008,
  14.1962769580769, 16.4055643066471, 77.5470624408273,
  14.7340227651054, 17.2470566225879, 77.4949075826086,
  13.6713373649259, 16.3976363657081, 78.3981650029753,
  13.3696064091047, 24.7331685281993, 62.5776184118939,
  14.1463022633593, 24.1419444931629, 62.3603681175812,
  13.0710758451053, 25.2088467990027, 61.7502069755192,
  18.576715941939, 9.33947253279174, 74.9237811756574,
  17.7556884791953, 9.85027595409479, 75.1787199334123,
  19.3406511565373, 9.97382636939307, 74.8054671955624,
  29.3008976004289, 14.0579052684162, 71.8487083729971,
  29.4423193890801, 13.7089825717439, 72.7751277323812,
  30.1670715859008, 14.4019364450687, 71.4862374412208,
  8.31872421249857, 27.7362210419092, 77.4525996295346,
  8.86839643317497, 26.9121691115385, 77.5897085857303,
  8.48404094994157, 28.0983816952105, 76.5352610674313,
  12.0345204049754, 15.6015686019111, 68.5153850102348,
  11.6984350871035, 15.0223058741512, 67.7727536404832,
  13.0218422365811, 15.7277139078088, 68.4190368777429,
  9.44243596224632, 11.6127000158523, 73.3901086318424,
  10.1588626740825, 11.916419036695, 72.7620262145228,
  8.99011620119179, 10.8040838662436, 73.0138816307491,
  28.4277916149106, 9.33800964989966, 78.8561579130162,
  27.7266984260213, 10.0508054559725, 78.8759184630587,
  28.3881119035584, 8.80784355856764, 79.7031227506032,
  14.9681872226011, 27.2524027876738, 82.1348790587659,
  15.4636960580229, 27.9804225745934, 81.6611088783278,
  14.1695935834765, 26.9866424235009, 81.5948608846417,
  12.2997579474137, 22.9035257389187, 73.3256789176362,
  12.8517224323643, 23.6910095314965, 73.0514445584093,
  11.7818048241576, 22.5690888613853, 72.5383565331869,
  6.86703481828821, 30.4689960114568, 59.8312086697498,
  7.80644843810626, 30.6334895404813, 60.1319476426306,
  6.40270978366066, 29.8818952450889, 60.4943187302589,
  3.32974051688506, 16.3169445769214, 66.7219748129628,
  3.95161324278419, 16.9102765764322, 66.2108667508671,
  3.11132601682532, 15.5105898779642, 66.1723502086797,
  10.6991469204974, 28.6168313144337, 83.8950618690908,
  10.6382452143707, 27.8016570507903, 83.3190567457766,
  10.2676735997807, 28.4338029158591, 84.7784255421185,
  18.9194350493739, 5.51211079043369, 66.2922112531059,
  19.9072339793318, 5.3582736080308, 66.3164474921815,
  18.540690842543, 5.39160081164689, 67.2098332726787,
  0.288210951246582, 2.84806923012752, 80.4236049727788,
  1.16455056109609, 2.69679189598572, 79.9662822679152,
  0.110562064462795, 3.83010321924842, 80.4872455041702,
  29.9842625024773, 15.5949643430639, 136.531782711876,
  29.3087827815309, 15.9747547084331, 136.773377621612,
  30.4331699328113, 15.5335446865544, 137.242140679271 ;

 velocities =
  -0.288258918958739, -0.0464757846202114, 0.309898594140005,
  -1.14126066542848, 0.136889613016801, 0.877358553021291,
  0.889648289021101, -0.128659109413144, -0.340988003387117,
  0.29095277052806, -0.121598980225798, 0.00781701565517309,
  0.111914091591883, -0.68577485140531, 0.281320962781623,
  0.050986017492211, 0.289902755264464, 0.109412916256855,
  -0.207717264495987, 0.217271141981879, 0.118045796372698,
  -0.702456126770042, -0.0425853080602091, -0.311184400699718,
  -0.411402279893897, 0.120738909058163, -0.0649355648292115,
  -0.147262570112925, -0.127364197866654, 0.0174020455144699,
  -0.0954313437465213, 0.317474001861963, 0.941217449358473,
  0.191869012350627, -0.604910464231653, 0.211270586973049,
  0.142034630565325, -0.0213885307871284, 0.175797920049009,
  0.0745881748867806, 0.117825914417918, 0.14820417585897,
  0.099415781022773, -0.0677062687905834, -0.00869741303930559,
  -0.195687224065716, 0.162271927774414, 0.0676033622836276,
  -0.332510212021113, 0.51383558357654, 0.761778954226458,
  0.17290027124812, -0.562951059444726, -1.38480505248441,
  0.025967413970105, 0.215459937423776, -0.307418361785855,
  -0.932843038379497, 0.489397009188454, -0.302692625326757,
  -0.0205445544744942, -0.652981455885074, -1.07716750039851,
  0.182652755124196, -0.0598060817655348, -0.0600669551077249,
  0.0495739389043515, -0.638149895948025, -0.345611732649458,
  -0.0230099997963264, -0.81615672927473, -0.413860248026064,
  0.159697103089859, -0.249762482369288, -0.280393523329485,
  0.276162896603028, -0.696699192360567, -0.0432190286352448,
  0.871473188367165, -0.200827230210862, -0.0427839048855081,
  0.110073767531674, -0.218435891800166, -0.282453698904204,
  0.652360574299086, -0.500184721076765, 0.396083036676587,
  0.279126111035768, -0.923061912138253, -1.05817360801991,
  -0.0698414348017167, 0.129122202269397, 0.228864682681513,
  -0.0797516801334151, 0.496570589407534, -0.819633717118867,
  -0.43190527454942, 0.753437469765031, -0.0222804556068844,
  0.0236033903264663, 0.0525034061339117, -0.171722650133626,
  -0.187337807796625, -0.370367925530435, 0.00586673014322748,
  -0.528439307061931, -0.497375209175789, -0.128526164911901,
  -0.10270506998053, 0.0206797155327327, -0.117844743712358,
  0.303585277608364, 0.537087446893001, -0.00781571597715667,
  0.431683479894554, 0.241717131896796, -0.697760976343968,
  0.0547035545928879, -0.281179260611942, 0.212650707835293,
  0.0736006716780503, -0.024819423809474, 0.0181128533099389,
  0.0367451546293814, 0.806109359504825, -1.12559266123626,
  -0.260819333013082, -0.174451065644216, 0.182115212531167,
  0.376069226050233, 0.114161439811242, -0.283141983832319,
  -0.0530756364742449, -0.683360838061527, -0.269195436523291,
  0.140585086485305, -0.0355571940065025, 0.364292852611372,
  -0.106381477117121, -0.210701290712518, 0.00142417290076508,
  0.077255733037837, -0.276195571735646, -0.0413813180100973,
  0.185602616162736, 0.198744236688188, 0.0348076217243044,
  0.940810260895477, 0.210443468515969, 0.391653453192079,
  0.40145445868709, 0.19439071036839, 0.141195563000751,
  0.076835016997977, 0.0910181835493285, -0.253087439909079,
  0.0754302245324354, -0.0727072945497582, -0.46590085923767,
  1.88220069010158, 0.195750928323012, 0.520283036194411,
  0.13845684847494, 0.324259735803958, -0.0137389557012224,
  -0.0396765657516758, 1.42224410349819, 0.777857422148036,
  -0.691273825033636, -0.369885899463474, -0.787594973866567,
  0.185969377643033, 0.0530349445010502, -0.233191623673194,
  -0.170154309994166, -0.551401710802434, 0.487648165146645,
  0.0851533800832843, 0.720480748254398, -0.738995663824711,
  -0.265357363511402, -0.01309620717001, 0.0652502213408837,
  0.63090764121555, -0.420557220816579, 0.266114597992155,
  1.10839638785501, 0.130954465368142, -0.0310729173991101,
  -0.0639512169064705, -0.263845739518765, 0.205325603283057,
  0.457164380792444, 0.146703635640445, 0.0845042077427073,
  0.0121246509301236, 0.169601666881395, 0.585808453962173,
  0.0136674314529313, -0.174643451554976, 0.122087155292295,
  -0.610369849325508, 0.0840398499725352, -0.44224824818083,
  1.04802423996015, 0.464840556898963, -0.244118020667926,
  0.15057316728822, -0.0105660543645467, -0.118831913887919,
  0.451267677522545, 0.203404878557359, 0.229761525917512,
  -0.11716185439704, 0.354503449650847, -0.273533642574485,
  0.0385857239857551, -0.143474243545149, 0.194551860727783,
  -0.218844391960137, 0.938467085838782, -0.91090749915162,
  0.193488532742659, -0.31192166625529, 0.404857200249924,
  0.253166257767113, 0.129804107189477, -0.232770062172323,
  0.67902056307923, -0.22948129170929, -0.0920556856262566,
  0.142965926391506, 0.43398688679998, -0.659743940726247,
  -0.151842292207405, -0.155549654571274, -0.106322401110458,
  0.706890811481924, -0.41583137396448, -0.0417958866939524,
  0.775354431347617, -0.438473477703464, -0.0251330862190588,
  -0.0564388357177319, 0.14979624975974, 0.0844868998223913,
  0.346334050977327, 0.301313745260838, 0.649346141765258,
  0.431219496510322, 0.467607033329838, -0.176124943992077,
  -0.00370705547149974, -0.0106928603052042, -0.281094339911036,
  -0.0632224484229247, 0.257373501802724, 0.594420728131647,
  0.131877665122087, -0.0280990174661384, -0.5611524043934,
  -0.145898992384636, -0.340243330549967, -0.180140327150867,
  -0.861544018691281, -1.18462602568541, -0.000156810956061295,
  0.321647148360482, 1.09518636592218, -0.957210602439821,
  -0.157119577143249, 0.489530889633335, 0.110233348036209,
  -0.232200079002809, 0.261612047817416, 0.449386270870639,
  0.0334677466934433, 1.53109045923324, 1.14996563480797,
  -0.106532250789209, -0.24846045560939, -0.0344245591525008,
  1.37574990788856, -0.594192233157957, -0.484667996249869,
  0.516534041574052, 0.174999706959934, -0.400254689585401,
  -0.131247052137794, -0.225851733201461, -0.0221302377013156,
  0.582510717666299, 0.586078778128516, -1.18401902796314,
  0.10542296695966, 0.165178043617303, -0.968076742220326,
  0.0596312559677408, -0.0486287119508085, -0.159086722445013,
  -0.0227250106392426, -0.192923714034306, -0.61112351009666,
  0.531434269832322, -0.378870187170379, 0.0442329617484065,
  -0.318692851487098, -0.270043554934513, 0.0146187343719743,
  0.657955760105923, -0.62733380560062, -0.023406848338784,
  0.503466314809626, -0.553056853400517, -0.0142267836514838,
  0.151072714879671, -0.139096587183337, -0.0700667651376435,
  0.208897154752068, -0.204092356372625, 0.267399127097113,
  0.281525746336, 0.0894990659525515, 0.203058953960893,
  -0.0471514616924823, 0.0455115833291541, -0.0888419321873047,
  -0.00457027474379722, 0.854732723798978, 0.197607617785358,
  -0.410176353101024, -1.06558857153395, -0.0960153547129882,
  0.130640976346638, -0.129067746343602, 0.073583716278984,
  0.0496040062918948, -0.22267212365932, -0.209950530561787,
  0.267973398909964, 0.0423221601378967, 0.0587600745813334,
  -0.152086273205074, 0.0313242386377557, -0.132051318198362,
  0.792190575118522, 0.00892975309253992, 0.00398006590705171,
  0.262531806273922, 0.424701508558577, 0.137023242252629,
  -0.350949814893987, 0.198445012282403, -0.0776370793503703,
  -0.736807881843256, 0.28623491832506, 0.82019891332237,
  -0.774288653636973, -0.188433141905728, 0.518227849539455,
  0.0991239141030151, -0.00361384389759939, 0.282375891705415,
  0.113057604670282, -0.989586567924898, -0.281434860151195,
  1.15769609450979, 0.254058624420527, -0.0862986243115222,
  -0.105355117092095, 0.115389010996095, -0.305809853585227,
  0.888567207064556, -0.0651014244341179, 0.588038338600599,
  -0.102472629504733, 0.969495277380978, -0.129763617633338,
  -0.234174085196851, 0.160196389586403, 0.10317518227844,
  -0.404836655995546, 0.00599160084319409, -0.231391384227675,
  0.158945050879559, 0.397893142706551, 0.107527276477409,
  0.419607166527112, -0.00859684956152366, 0.416300733950345,
  -0.429623242119729, -0.140783642598772, 0.0786862938327756,
  -0.761723209873073, -0.155882858740721, 0.0516215382231428,
  0.0992748182965588, 0.151523424095654, 0.362636795618951,
  -0.292533677444276, 0.601144989731425, 0.562325410947757,
  0.264470933051756, 0.0896131277529322, 0.265318052902586,
  0.148957893075978, -0.176824529041887, -0.0294332760419921,
  -0.620851501699761, 0.0932957688486337, -0.332496140617227,
  0.234412379789785, -0.103891282218437, 0.350660146699398,
  -0.0573279801763814, 0.212503784729644, 0.504175079000992,
  -1.10224066965622, 0.124558558400531, -0.827884478941723,
  -1.15996416731471, -0.0074175716541191, 0.231874348836485,
  0.213561116803051, 0.176683761632773, 0.242786650152856,
  0.0728512651470099, 0.524575392428188, -0.0602996415044297,
  0.185315455024358, 0.16263665954147, -0.349375764357728,
  -0.11930474475603, 0.401016267602, -0.114569310539074,
  -0.314518110875313, -0.0268303088244554, -0.480432169395732,
  0.213406791225785, 0.67409886458773, -0.235298481679863,
  0.0811489097364827, 0.162328396160729, -0.157646541488832,
  0.0193863874300564, -1.25521722031524, -0.201117313711166,
  0.995755275556308, 0.367551292734466, 0.608423713203723,
  0.0728455418354761, -0.224664330333633, -0.0918135723321132,
  -0.177298060955239, 0.216077289169686, -0.346091195696718,
  -1.51394530688487, -0.0419705032260555, -0.836705677115679,
  -0.170007621518867, -0.0800400247314791, -0.0988235446949705,
  -0.462619830698482, -1.17176342755202, 0.442163959474774,
  0.101002475185018, 0.355254949282777, -0.259450783068543,
  0.100258442040431, 0.0019097198626025, 0.201581263102155,
  0.513688452596184, -0.636835200499204, -0.130033998112712,
  -0.665438786997717, 0.0380978377609156, -0.0751842311701411,
  -0.0227355411438078, 0.00653209385926725, -0.0691188575576798,
  0.475214570920024, -1.13540128261153, 0.400354390361133,
  -0.294039828887521, 1.03922200045371, -0.580634780119168,
  -0.0862952031424733, 0.0209321077442984, -0.34745896486476,
  -0.121804767447364, 1.0497801665094, 0.121258634363742,
  0.524118743243235, -0.549450147704993, -0.225631155283899,
  0.231278497136979, 0.0414893215748298, -0.148613057963537,
  0.34172707555109, 0.511812777020914, 0.549060107180386,
  0.438922748925063, 0.208784451300456, 1.17228911198787,
  0.22555373083152, -0.0381866893613945, -0.16701492217435,
  -0.0609182640293406, 0.397651941783735, -0.707276533368903,
  0.59045818622945, -0.746132040539624, -0.431431468370588,
  -0.131645905646705, -0.065278979045236, -0.31311247771162,
  -0.35262137324626, -0.193433600236368, -0.336055683122003,
  0.201353546283115, -0.0844912186665519, -0.474614885889875,
  0.0802455679857827, 0.0442704773163313, -0.0220916542956472,
  0.225130835624132, 0.147292304582755, -0.370647746704906,
  -0.205696607846851, 0.162143399256304, 0.187053688453618,
  0.239940040992457, 0.171153329457676, -0.021012448013134,
  0.68654403626534, -0.437699071001338, -0.669934935007159,
  -1.22583833134622, -0.22477872179128, -0.379677241736894,
  -0.4220050766227, 0.0918474143445507, 0.21144286290617,
  0.180796576514287, 0.207031765980837, 0.678285691879861,
  0.352995393139706, 0.994751797952279, -0.27587801122296,
  -0.299283242143206, -0.0504241701790083, -0.013672528973121,
  -0.185994615022801, -0.138104990912195, -0.459918776511811,
  -0.206992288207593, -0.190690913074393, 0.106056806802489,
  0.211140635638508, -0.0548427310518329, -0.34560478614642,
  0.257755859366418, -0.168560129065061, -0.558301706260162,
  1.25705953020371, 0.704623296700123, 0.0415653878386203,
  0.119297392158106, 0.0499395129528446, 0.273267455438011,
  0.143188126719228, -0.684346141606498, 0.220707950182662,
  0.601899703726388, 0.266048253879062, 0.785329186298136,
  0.177120553171771, 0.224156731277041, -0.35708999123685,
  0.0468971826553068, -0.328967140308411, 0.0485615921053763,
  0.0498095956659973, 0.806569912500668, -0.013695129980376,
  0.26831267420513, 0.0654425921452292, -0.0708736904677073,
  0.132403262731337, 0.121507883281443, -0.553133443195747,
  0.781589129789984, -0.371062388027123, 0.373045402379234,
  0.222143646711347, -0.009723474866427, 0.378688962686707,
  0.722211840942252, 1.1110743526128, -0.168594162827556,
  -0.695009217049958, -0.846779800181097, 0.951371715673216,
  -0.168533900119171, -0.193985318637625, -0.174865262090693,
  -1.16326938746647, 0.0506573566579289, 0.0794530546118311,
  0.851258640863181, 0.0264418064220077, 0.299267427333792,
  0.0536135422709361, 0.0911652477339779, 0.240103232748727,
  0.0277260345626171, 0.229466710084135, 0.276109804456157,
  0.682834773650667, 0.616062840122916, -0.707011682042351,
  0.0709159766595508, -0.0308960731705039, 0.0835329338188096,
  0.0850429752712908, -0.714459447399135, 0.684524146938789,
  -0.0529959548865148, 1.18061272634899, -0.567135586158487,
  -0.216855297529962, -0.173735734906765, -0.132460912213255,
  0.236567752270882, 0.158514072118127, -0.278862829563683,
  0.0989503989045104, 0.287142167703973, -0.244503630768348,
  0.103936827346713, -0.242140661862201, 0.149639262349483,
  0.312519615205179, -0.0927144418208569, 1.01172326818634,
  -0.314167169225732, -0.254080777275226, -0.98828316173095,
  0.106159995687396, 0.0468152245539133, 0.224748886692853,
  0.187189793202448, 0.0076331981367108, 0.779554374528872,
  0.193091423810344, 0.580489642662765, 0.0190993018971334,
  0.0235626337936209, 0.21020562490307, 0.0726549004612771,
  0.375708273545945, -1.31509028458113, -0.24128849793512,
  0.163458926960176, 0.80947038267814, 0.112010409867045,
  -0.014571300106089, 0.367577098250033, 0.208058978251158,
  0.916408140873248, 0.192450175684646, 0.598586940731359,
  -0.325351742793835, -0.0997517284322876, 0.629842718358898,
  -0.168764377369211, 0.167235476723829, 0.0834058479263984,
  -0.452975109663432, -0.533014252877721, -1.40943202675246,
  -0.584723795711649, -0.939917515727906, 0.596402345919479,
  0.13664147512268, 0.0869818438448241, -0.0915751554900498,
  -0.542997227752864, 1.03107439290745, -0.575368560807159,
  1.16722681148566, -0.209364395165722, -0.751330014074511,
  0.0607283580287494, -0.0641197011501244, 0.228142798933374,
  0.734032776580181, 0.641062312698205, -0.364908895067551,
  0.596508134758197, 0.857170760678885, -0.106510857110084,
  0.161131354835903, 0.453884138596452, 0.336937663660309,
  0.11200654826875, 0.707152359921084, 0.812327047328526,
  0.624758375635803, 0.127204744507736, -0.205508530534893,
  0.0119176212756483, -0.187562891896342, -0.0820791180456568,
  -0.219045616897303, -0.120507490943029, 0.372054964962479,
  0.116762281163418, -0.0512582298443732, -0.161357113023223,
  -0.209875076388315, -0.154497485637194, 0.47774130730727,
  -0.767315163832267, 0.177344453546396, -0.246290868657383,
  0.499083828690404, -1.41109546902718, -0.568314587880269,
  0.266095224826577, -0.165357064100599, 0.0977422901958189,
  -0.0421502242024275, -0.657785182024309, -0.113736210496585,
  0.831518135145842, -0.192451519645575, -0.0744169450729985,
  0.17342354151146, 0.0421324037971495, -0.0275677770912183,
  0.127149488900395, -0.367746161415629, 0.0291101511816055,
  -0.502366651454818, 0.552290604965675, -0.728042239737218,
  -0.320142247308928, -0.242231676134124, -0.125454065075445,
  -0.954641051699605, -0.467201625318725, -0.276667198780926,
  -0.594302297020747, 0.498866832368995, 0.752443889571556,
  0.0993078995349185, -0.258575395960403, 0.123994249207789,
  0.57333203071459, -0.244811469371323, -0.453644205614677,
  0.0295695888645171, -0.391970795399498, 1.04995048511661,
  0.0719175300239694, 0.0928213062390161, -0.0234277638782275,
  -0.313687915044863, 0.526031711757073, 0.554072861412578,
  -0.253146012452011, -0.655448635164179, -0.0593664728630183,
  0.0244165623033703, -0.296974020351947, -0.209985089958474,
  -0.462416227840082, -0.0371242705133566, -1.28442170404857,
  0.208085821822593, -0.398568938366468, 0.150930256438767,
  -0.33800432156584, 0.349179940776081, 0.394327629472261,
  -0.416902341639837, 0.582953317969973, 0.669667479569097,
  -0.526763023952002, 0.0983489575585267, 0.45629054411122,
  0.116794058337189, -0.215441746766767, -0.104165663248286,
  -0.445317567182456, -0.0733428487014696, -0.894934648076645,
  -0.359480293283306, -0.192079351999137, -0.267194715165097,
  -0.136880539691098, -0.277909262678087, 0.024452587203221,
  -0.628015566119693, -0.523507613102635, -0.0170871262961646,
  0.771330644583694, 0.22729851566276, -0.482444724499121,
  -0.307005909439731, -0.19716297115204, -0.250540515080372,
  -0.664480099445993, -0.0551378450976168, -0.330417003368103,
  0.426048780946084, -0.495082640693599, -0.0809910042430923,
  -0.214069979149265, -0.0782200014237289, -0.0065022937431078,
  -0.990116483400835, -0.232743035640215, 0.790911114646288,
  -0.0214743240011671, -0.182857690271502, 0.830478320707883,
  0.0827579337815852, 0.234639889699401, -0.376574381345542,
  -0.801710541306895, 0.791675030724926, 0.170118280052606,
  -0.0988424268636203, -0.406220369431293, -0.0948960630336845,
  -0.0576701676909147, -0.235342416861459, -0.0749689788334116,
  -0.122083392598388, -0.790947265565956, -0.939387585330225,
  0.976821502213171, -0.812873498898122, -0.244581818687433,
  -0.120319217648587, 0.0469364491087813, 0.00381863011290764,
  -0.31703098324753, -0.248677570241635, -0.118421502256657,
  0.118638927732331, 0.252288562849602, -0.260729368504185,
  0.0659055208003713, -0.0350718575575834, 0.212652532484028,
  0.42489324704185, 0.307492084691905, -1.50209303233998,
  1.2127543734494, -1.32489062195442, 0.700415779978496,
  -0.0621068308444338, 0.0284534396533834, 0.00592561659668011,
  -0.312683722395071, 0.270891377924262, 0.810607012931313,
  -0.41109059762467, -0.0101697708848905, -0.139880943760461,
  -0.125778241084266, 0.11238439453398, -0.300383500208302,
  1.35392167344767, -0.603651262219056, 0.405848036166001,
  0.460448113953503, -1.37315734675873, 0.635197672844677,
  -0.038841995749933, 0.0593969276329553, 0.00606241309438166,
  0.117882271182047, -0.308836102529681, 0.311909192176311,
  0.226167352781057, 0.178729501101958, 0.179357679936094,
  -0.00876474071197482, -0.0833513640843155, 0.0668983700958244,
  0.321066143854823, -0.198345292535823, 0.0170707370185059,
  0.0692601502171447, -0.153149749543392, -0.510116696187786,
  0.249425566957409, 0.281152867272021, 0.00862114108212074,
  0.0818450765670127, 0.968479931116377, 0.840883199640353,
  -0.921279689278693, 0.120363502084821, -0.387327050555928,
  -0.223405785293506, -0.0487693287448368, 0.299496094231056,
  0.471505725881426, -0.211576408297608, -0.161062748235809,
  0.626302069324935, 0.440565113093408, -0.161376236074718,
  0.140733333068298, 0.00796082178896303, 0.213161034035582,
  1.02855050238316, 0.522036597827463, 0.095530986900555,
  -0.672276468369366, 0.716181366571483, 0.309669787082237,
  -0.0462824342700047, -0.210851630006958, -0.326938981428275,
  -0.0852142735381626, 0.0463890898546214, -0.618074623662868,
  -0.0840970024236439, 1.01127408311093, 1.12114660046545,
  -0.0139317179226928, -0.0799210299511606, -0.18714309406432,
  1.10829460888124, -0.0361423087942488, 0.47994681364579,
  0.140641915971988, 0.151916459496017, -0.375005837036986,
  0.197073779660486, 0.131269445676297, -0.102860998684282,
  -0.12526704039334, 0.465387429078856, 0.492178916832735,
  0.547811210102982, 0.0223774486341666, -0.251486711274648,
  -0.0558446842367906, -0.0456303681282671, -0.114651648257694,
  -0.15321193091232, 0.136670981654882, -0.108172483363215,
  -0.110897579461041, -0.210898013044557, -0.383519690661653,
  -0.21888835757601, -0.0707636703844709, 0.289310155307303,
  0.347847377691016, 0.683498279372246, 0.130429397358494,
  0.218627110189908, -0.562485054471796, -0.514607599285295,
  0.179906623184017, 0.0776775493842997, -0.0043982433962986,
  -0.0517778046181051, 0.608841576227528, 0.416426954394062,
  -0.366903453165203, -0.182899304397775, -0.379876636004731,
  -0.0859701490925265, 0.154662179505167, -0.0846725108071661,
  0.373974204262929, -0.44717860127321, -0.682435985512079,
  0.278902455561742, -0.282000816468688, -0.531751574314367,
  -0.116194450432103, -0.331053404481893, -0.28686290168248,
  0.081349731256194, 0.12805397465955, -0.381061986925894,
  -0.152869428226903, -0.406474572779818, 0.388227533244273,
  -0.0909435862629968, -0.129687097328702, -0.108458399960417,
  -0.0977498568964568, -0.00243054974841911, -0.1674307662548,
  -0.0389851789623176, -0.148631894794576, 0.0115116895512045,
  0.0322846457127568, -0.0862525528038172, -0.187783002457087,
  -0.615397483852399, 0.265469995237538, 0.183436521513078,
  -0.467482589193808, -0.426241342711134, 0.402746819100381,
  0.0728803277055458, 0.0736649167158579, -0.233636251323333,
  0.526568572503843, -0.509411380313638, -0.616077625139756,
  -1.11929576012586, 0.687682852593903, 0.634030614509125,
  0.036481040728258, 0.11004371068764, -0.135310531610968,
  -0.460736098578216, 0.889663949000414, 0.752033528907971,
  -1.18647222734219, 0.383738245994587, 0.319779439738951,
  0.115795195821732, -0.283503533575113, -0.145838355812407,
  0.0523872995251008, 0.0231453606002685, -0.327112428419193,
  0.192320318513865, -0.65385783881128, 0.0731449447813894,
  -0.0160245942344052, 0.11224390975786, 0.0259517685966919,
  0.955938650470589, 0.430323383379997, 0.379418574213577,
  -0.437123602383807, 0.945327123505469, -0.432332960573596,
  0.0332075644780744, 0.206607139133576, -0.291128690401183,
  0.471172791800112, -0.0175093819923599, -0.437969179436112,
  0.303018359789946, 0.102826940789811, -0.277117322543563,
  -0.0122990194751698, 0.138833323359754, -0.151433322567308,
  -0.0387805720997369, -0.323128634712118, 0.481735696361884,
  0.63795230371765, -0.976236232174529, 0.232168260281307,
  0.250859082066813, 0.153404167267359, 0.117815056090888,
  -0.0448959275897231, 0.670019587928286, -0.338719881713762,
  0.452956997713294, 0.216236878539592, 0.0833730209614274,
  0.030076204915108, 0.273019053434387, -0.195699167012177,
  -0.685456314281502, -0.257240767356133, -0.00255003982409283,
  0.789569315466827, 1.20106717443067, -0.151421916738008,
  -0.288609736754911, 0.0513319181751561, 0.0926923372822603,
  -0.413171447654687, -1.11099138087828, 0.685379701358635,
  -0.0211667417113301, 0.22429284202215, 0.588620020180625,
  -0.0245050716589823, -0.177825784011878, 0.157088231721019,
  -0.398096299377156, 0.354161235464821, 0.856381264241861,
  -0.408047231258473, -1.07162551920273, -0.61492302820023,
  -0.229971445172852, 0.184549804325168, 0.0442576619646399,
  -0.220838330669275, -0.604291764011364, 0.0199959995078246,
  -0.154866622977069, 0.384672028729983, 0.126906492306713,
  0.0503410583994568, -0.0837175104041625, 0.107605099903876,
  -0.262550556891082, 0.0813124173486909, 0.363111960335281,
  0.083519047073882, 0.0158359517229128, -0.114224054892671,
  -0.0323839972676331, 0.227014436274452, 0.223947508103585,
  -0.596168832943425, 0.961803597494142, 0.486573923251674,
  0.428445857052013, -0.560044876862925, 0.265798614024083,
  -0.0533363723887683, 0.299781348588186, 0.230964193228188,
  -0.131248726043481, 0.368538456857474, -0.831371715893096,
  -0.242345186842917, 0.0637203757722294, -1.29763466836752,
  -0.168310360063035, -0.286184895395933, 0.235772639415584,
  0.0576044234423242, -0.434994071211063, -0.58211511942652,
  -0.0415839160335849, 0.381878125520238, 1.26684399897285,
  0.21388989049625, 0.0135369092033, -0.291242060285086,
  0.33159611728269, 1.09056001755317, -0.901972604915913,
  0.216402260697991, 0.601892445288055, 0.291014906448196,
  -0.385070542066949, -0.00096098737639104, 0.0834674344787206,
  -0.207047505558782, 0.0784814580664037, 0.644970354315033,
  -0.313313016679783, -0.248836521110605, 0.113319278023064,
  -0.16106038860215, -0.027015955602712, 0.280883171942425,
  -0.372238751956262, -0.0980785754045319, 0.227165270009894,
  -0.571627895227281, -0.350045135387101, -0.0386282504951013,
  0.090063520297507, -0.044735271007381, -0.0146704530231508,
  0.424681605929501, 0.552563516665747, 0.222669717879723,
  -0.460039020497817, -0.399662545798017, -0.453944029451388,
  -0.100186961741514, 0.0934440028481948, 0.0472453780361975,
  -0.535386762633772, 0.353046674149531, 0.761155439094279,
  0.0347738131717256, 0.406802372995601, 0.542404771109918,
  0.146571367681313, -0.253073292723318, 0.161004469772117,
  0.124664884285003, -0.503790423160767, -0.0555895179931331,
  0.184840409770088, -0.0225832157532005, 0.211869043983182,
  0.0358016903857546, 0.0767087145896558, -0.0595060671136234,
  0.201971630462569, 0.021611440327163, -1.11320099120558,
  -0.92705164247626, -0.314325621262482, 0.165541081437365,
  -0.206347051420201, 0.0889302571989347, 0.228243066926462,
  0.566877550853118, -0.161387489041196, -1.56507435743326,
  0.375262854603302, -0.642979294714183, -1.01631934590505,
  -0.29468267418101, -0.0751360411193483, -0.128598738925057,
  -0.193709510717799, 0.0624783649489287, 0.0849271495833923,
  0.213467395411191, -0.682364728658879, -0.0815149948912531,
  -0.0472200510384237, -0.130336195020737, 0.207098252272515,
  0.139397085510642, 0.0848703370708392, 0.34438114489007,
  -0.425713733658872, -0.157441208774325, -0.0845236770266885,
  -0.0028420891320382, 0.142662569760575, 0.0669584624981787,
  0.0696638872820661, -0.431010275996093, -0.0289207861989523,
  0.53668217817677, 0.697016198424314, -0.317676606642337,
  0.0456451452148749, 0.0611011121738533, 0.161265219026208,
  -0.630326155011763, 0.811482640156697, 0.234337495817305,
  0.894025739195213, 0.619320009244671, -0.455281042371212,
  0.29670140030787, 0.110570629190712, 0.0422214221608231,
  0.269444474974664, 0.703842629338606, -0.00809803484169211,
  -0.462840504332388, -0.460976722226374, 0.233798367604828,
  -0.341871957574501, 0.140546408109243, 0.339977124710119,
  -0.081639975295996, 0.156032006616736, 0.557243356746472,
  -0.304439646658127, -0.959253249588137, -0.860337542001383,
  -0.335818588344307, -0.147342314071709, 0.00639653947396196,
  0.0917451917044096, -0.446118479812005, -0.0172214206580038,
  -0.23849444154141, 0.315560082207083, -0.0347178494742454,
  -0.0564023106742137, 0.373572063617986, 0.389358529621289,
  -0.285560992803811, -0.20786859825812, 0.26956608438751,
  0.117473778448125, 0.0875584165663933, 0.966370082436245,
  -0.00197608015982122, 0.132129168870623, -0.0287046689172132,
  -0.801419156544139, -0.585492833721465, -0.0444296777679089,
  0.369607731259253, 0.631444696408322, 0.177658703608578,
  0.194036191474864, -0.218146279955038, -0.291293055225473,
  -0.406467176034629, -0.197587969525718, -0.312861940777202,
  -0.372917045712317, -0.0277466659964283, -0.146917599162637,
  -0.103742597791923, 0.347534982170792, 0.202700356647893,
  -0.465200939842678, -0.104986792401975, -1.13944631211785,
  -0.264064989865707, 0.0898179039049683, 0.110210059748807,
  0.232068544014319, 0.110190803621524, 0.407394523758322,
  -0.334537805145968, -0.226348408775872, 1.24158938834068,
  0.787818361505815, 0.140551024183973, -0.542815918275011,
  -0.0445500475954449, -0.294377363921237, -0.0821978551043439,
  0.793665032879286, 0.183554038589427, -0.287208210832699,
  -0.558408693461986, -0.0432815697999088, -0.154916703532649,
  0.022165706711548, 0.0471207995781507, -0.0187769616697588,
  -0.878802450265825, -0.917006054845234, 0.0789330310917168,
  -0.238678525644986, 0.457238046969272, -0.441508214176207,
  -0.0563778111447057, -0.0636094656038664, 0.131112242365866,
  0.570836454312683, 0.148713270914487, 0.696986732565809,
  0.160238193563929, -1.19198742828525, -0.599622161640274,
  0.125243569324465, 0.121522784420393, 0.429640065554805,
  0.334907925011282, 0.185492068662958, 0.474540704787798,
  -0.67825834660568, -0.125028773611659, 0.250889162728922,
  -0.0309943026098831, -0.0800147992401453, 0.367138288384173,
  0.637136361696317, -0.350120587132249, 0.231164532724548,
  0.436773087504934, -0.109417163297055, -0.310526242878083,
  0.420462522204868, 0.0368023742544813, -0.202878972905124,
  0.994270912972228, 1.135842187355, -0.988017899571402,
  -0.349480541868386, -0.186890173493519, 0.988176073886852,
  0.0912754754368985, 0.0299468604461558, 0.160306126184277,
  -0.134617786289474, -0.0532361333798229, 0.541368323648968,
  -0.184954163104866, -0.453411495096775, -0.505544859327681,
  0.166659401922507, -0.0459462577147131, -0.151941294279422,
  -0.168843461673128, 0.382382019714346, 0.257271208078001,
  0.24130360574166, -0.221558706741429, 0.095010682737076,
  0.126360670949096, 0.217534328411579, -0.00610852242767552,
  0.29983162288036, 0.669355082030965, 0.010544423639958,
  0.305463570873137, 0.0212010490298252, 0.415664782623394,
  -0.0563568869288598, 0.107281818007466, -0.339421517694724,
  0.246951232845517, 0.692799355138874, 0.35641812891156,
  0.169316795940881, -0.126425634850336, -0.105730344268425,
  -0.16717239351688, -0.24494626460904, -0.0690564880004628,
  -0.496337862405401, -0.192224543381322, 0.125773722163533,
  0.35059855837035, -0.424018022315131, -0.225775194855206,
  0.21480561548562, 0.0948316890239467, 0.148005606998981,
  0.663247248637344, 0.0404465241012647, -0.0866147984716148,
  0.32890703515085, 0.383079020755916, -0.397703541262535,
  -0.0545358010954589, -0.145794941330805, 0.189630191051908,
  0.178487397900613, -1.40155752047855, 0.0167741399319533,
  0.96054635889009, 0.0259143222205798, 0.512243838723317,
  -0.0653600186157382, 0.0844798355657834, 0.134946749752989,
  -0.953266221717205, -0.88461040237724, 0.53266721960224,
  -0.429329764051613, -0.901509465936691, -0.0654209602041986,
  -0.136970467133652, 0.0677286145737447, 0.156078304514759,
  0.251535007884273, -1.02790775620313, 1.57299396836204,
  0.858846584410778, -0.788051921503112, 0.589829738235179,
  0.12761322083965, 0.0761635103776581, -0.00571853821297213,
  -0.518329866743201, 0.223829943740321, -0.671716561605256,
  -0.521208206548916, 0.414653356157807, -0.273577744452081,
  -0.0783739961454807, 0.256585862459021, -0.0478160234414414,
  0.295265945999553, -0.506385606146509, 1.00425096952678,
  -0.181400079627503, 0.315541507987498, 0.179689374839474,
  -0.0573021668614421, 0.0633970060222729, -0.0121894673269645,
  -0.88715785660463, -0.273545855573211, -0.114082523654284,
  -0.406906925711861, -0.0716621381804749, -0.147320897402418,
  0.0102769679661627, -0.124624476392647, 0.155827486045628,
  0.526352612029298, -0.379533289044416, -0.0826849223219514,
  -0.700171904480336, 0.779619260491077, 0.0385610822330683,
  -0.203993110537815, -0.170652227692265, 0.158246533526938,
  0.537881736279767, -0.583297586428837, 0.804489525190462,
  0.225383506228851, -0.0262892983528343, 0.0711983005010117,
  -0.0244312702993582, -0.0790750248686315, -0.0852540767867003,
  -0.235310150315144, -0.968625843768, 0.21762676157332,
  0.258066547551795, -0.0570290753237481, 0.615051812879264,
  0.294049541990219, 0.268627712372605, 0.140734393458587,
  0.397536275944092, 0.565839123920322, -0.294011289876013,
  0.063973699420694, 0.424505836312459, -0.384656147147788,
  -0.0835322202945646, 0.266237188233782, 0.244760381138638,
  -0.402038118917001, 0.200034260297397, 0.115380865475899,
  -0.634037397918723, 0.786183286281465, 0.470941723884806,
  0.159761271618445, 0.0621205738447944, -0.0108443870421292,
  0.1581015936695, -0.707228956227306, -1.07172440732842,
  0.244827432041624, 0.410737284714043, 0.830121046526541,
  0.000594188982869377, -0.120238823094182, -0.0529712095370097,
  -0.280742020053443, -0.725437162866715, 0.374019194590946,
  -0.074210339847184, 0.219325058869524, 0.0662117692627195,
  0.0871333632151873, -0.261877339260972, 0.0823916506615497,
  0.586026585072436, -0.379561155116331, 0.133476261586937,
  -0.240243413036605, -0.444346793764705, 0.347627225163265,
  0.191852990277103, -0.178517867896503, 0.226001833590124,
  0.121783196400441, 1.01511362641454, 0.0305531552663225,
  -0.147064851136472, -1.25238030506507, 0.697716408564316,
  0.201560070631329, -0.128434969083479, -0.0893399473987531,
  0.298034185025648, -1.33384877073969, -0.484217736934228,
  1.20813683265137, 0.234182468292595, 0.256829372224088,
  -0.254711315565081, -0.259247666774645, 0.195240295819926,
  -0.514941688180837, 0.11146016004271, 0.577349685540512,
  -0.167140833143445, -0.380735171915738, 0.0254952071049746,
  0.0310636129550538, 0.253996660771051, -0.153428388570842,
  0.454628227382845, 0.671728805426184, -0.228434504319291,
  0.667465388410207, 0.353793463008133, 0.089387683071448,
  0.297512588022366, -0.308414788833874, 0.152572958556937,
  -0.717213233121036, -0.412991749857899, 0.590159181327719,
  -1.10069688207024, -0.601965074989488, 0.44256835616395,
  0.0520415723546095, -0.181957919534994, 0.085270098410338,
  -0.301696287830441, 0.809822130481441, -1.52004660887644,
  1.36676332765269, -1.19796633016921, -0.77454284868699,
  -0.0609164524929937, 0.217839533799622, 0.122263959536676,
  -0.0122930377648093, 0.14260282148727, -0.0569651747225739,
  -0.0190083919185253, 0.177870355407639, -0.11030821774677,
  -0.161957879170458, -0.00101800553448848, 0.12038309158717,
  -0.371748825623586, 0.0155677748887959, 0.417177248138358,
  0.132439104011209, -0.169570637490676, 0.658449777480192,
  0.129095809911509, 0.220972894665691, -0.112183569114034,
  0.00879152040172548, 1.43518943552167, 0.089667233364832,
  0.384916545672943, 0.130726564555637, -0.205549194356197,
  -0.105800671632814, -0.264430136280108, 0.0712923653900166,
  0.32819018577107, 0.116890668929911, -0.118781758097982,
  -0.392632037328316, 0.0511008285083223, 0.303818014900493,
  -0.103661638196558, 0.0696091877017708, -0.00571933849702963,
  -0.639419127880551, -0.124002305680706, -0.346474780608269,
  -0.177074862714275, 0.738522156989123, 0.0670968467037101,
  0.256202710645238, -0.156257097827568, 0.143044863477951,
  -0.254256163821589, 0.00319629669579863, 0.198573913442249,
  0.186670365514883, -0.214166661605152, 0.475528622190317,
  0.0296143598005128, 0.501210313912377, -0.081503666680801,
  0.291486587472493, 0.322216618464907, -0.739026590503838,
  -0.0614732740047315, 0.314819209404806, -0.27410403503763,
  -0.00767714269656797, 0.00205056673040339, -0.244873504434512,
  -0.101357360516016, -0.612041433006607, 1.53186498702806,
  0.493059462916085, 0.47368191463727, 1.72421271368637,
  -0.248564228755039, 0.0321424285966808, 0.238534188275053,
  0.352119152305872, 0.0700212556108845, 0.00782236935899736,
  -0.0557995276089579, -0.0358546507929705, -0.221281501834137,
  -0.131469667815429, 0.0876275644661409, -0.148274933916641,
  0.123746786848849, 1.48998538857607, 0.328736118654978,
  0.760132937147987, -0.480415519918226, -1.05905664033515,
  -0.131957632645735, 0.0137521337830264, 0.0676056718966244,
  -0.359119496251228, -0.057335293433755, -0.588215271158473,
  -0.0676304771331931, 0.148152505693347, 0.274576321817238,
  -0.0648656786606246, 0.0893131044723815, -0.0553870942621659,
  -0.219142979626866, -0.162146780466921, -0.172290840898734,
  0.754966816434032, 0.597157124974261, 0.750365575334825,
  0.12442929399905, -0.0484055863444716, -0.41090827037624,
  0.142714370781963, 0.47062475057551, 0.064297676970574,
  0.00154170186989073, -0.0948575834138029, -0.365117305681894,
  0.20188967534453, 0.17293806061351, -0.174386591458894,
  0.839770239194151, -0.404851953367715, -0.816846888419881,
  0.677967078105284, 0.100741803768119, 0.644994807488184,
  0.148594493171453, 0.172739030535624, 0.223190055473968,
  0.180788727592275, 0.0505576480910309, -0.162310347711767,
  0.288949323673479, 0.0362957464899656, 0.603212258289277,
  -0.0189751566936053, -0.0468345732623875, 0.213037142651605,
  0.940494907446807, 0.0821337737594474, 0.138383493021915,
  0.536845604997785, 0.583923996218115, -0.938506404258271,
  0.069899901360832, 0.0982829139132626, 0.097141656489165,
  -0.0899629517182028, 0.378330938988032, 0.252582951013802,
  1.25565053001818, -0.0645377349297121, -0.081483259628735,
  0.136348820123752, -0.123478759182892, 0.245542086968176,
  0.244721264494528, -0.139378118789469, -0.0803186532888004,
  -0.0126381895352835, -0.258910155583625, 0.322464444884952,
  0.360731965003953, -0.0654344801484165, -0.107387188224703,
  -0.265032601749, -0.250911692334708, -1.13246242426965,
  1.03863632732309, -0.964043726678332, 0.0858531216583127,
  0.106858584582083, -0.0688257494234087, -0.476996535885832,
  -0.360104296167033, 0.165636253798929, -0.909099934513833,
  0.446845358382832, -0.412736178609121, 1.22801863445149,
  0.213198856877764, -0.120989868065821, -0.0479347319478084,
  -0.324796826551033, -0.577952410036187, 0.285317471552476,
  0.105951545944223, 0.746955868839002, 0.933365938142564,
  0.0074183430385285, -0.15066089408922, -0.0237780808280482,
  -0.513071281633835, 0.122121382047177, -0.139731846776266,
  0.659619675275301, -0.0022309193939465, 1.82201493686731,
  0.0114887067671319, 0.0447693589043393, 0.333285821197715,
  -0.186371187533035, 0.577192927759743, 0.171797230844521,
  0.0771296950948768, 0.369263961983061, 0.537686300399615,
  -0.288012949565104, -0.126426520657302, 0.112602389672767,
  -1.17623506493774, -1.34524195079669, -0.0304055590081325,
  -0.676723277119017, -0.234745548534668, -0.311189438885746,
  0.0407201322567075, 0.15340620466763, -0.162327829102815,
  0.275468716223764, 0.477017270099841, -0.243295338563775,
  0.010509103507534, -0.0238243936494226, 0.010888100997087,
  -0.137247144390297, 0.0045364914109263, 0.536354124753304,
  -0.0232355912445724, 0.134149571662243, 0.55862269487859,
  -0.100115209988177, 0.0407874266738144, 0.520575264643645,
  -0.270582619845867, -0.163739046852085, 0.174990216256244,
  -0.287007524606302, 0.112147090561044, 0.35521328026977,
  0.0714883868889922, 0.0651187008288112, 0.532663052160195,
  -0.154750007945296, 0.219447241332829, -0.291618872855597,
  0.222686654411977, 0.507720515679312, 0.0283473220975967,
  0.0575328819415527, -0.0763289752017595, 0.289262718485652,
  0.152368747367139, 0.106988381589815, 0.167084545618761,
  -0.593050702736232, 0.904684172893416, 0.104194843355358,
  0.451609340899675, 0.0567642115725554, -1.22103349035402,
  0.18334441351973, -0.0396147410876857, -0.280851670257241,
  0.919387242248083, -0.160469386041232, -0.67058262318844,
  -1.01719588678383, 0.0578234012793226, -0.314099530714498,
  0.273068786572736, -0.0436689855441508, 0.104014686460497,
  -0.240508351188491, 0.315792539950048, 0.243557229838069,
  0.426577627972517, -0.0804519192950918, 0.672125626839491,
  -0.175437250704118, -0.0520757251490346, 0.0283985967052424,
  -0.0181828458339728, 0.670746152751812, -0.373507060623348,
  0.0704084091851157, -0.17438483283792, -0.377365271008198,
  -0.252512127611905, -0.0913387694626674, 0.124597510583458,
  -0.880022193525066, 0.556622396330144, -0.101208855162207,
  -0.00779335397000858, -0.0927712576145899, -0.176060765439949,
  -0.104048037526223, -0.0223217770844693, 0.186400591137842,
  -0.462564305748853, -0.323096934434407, 0.423120893050509,
  -0.514227582679822, 0.0150839633609827, 0.570440187658873,
  0.086326842057118, 0.0588743501661512, -0.00205446700664323,
  0.253956129879727, -0.532473737552955, -0.201126679978867,
  0.423994296235783, -0.0720472997488411, 0.124706012376337,
  -0.0716886439544052, 0.0747576648398886, 0.262444266237723,
  -0.0172819725749974, -0.291115830138644, 0.692272501822237,
  -0.082876280301252, 0.085319165105237, 0.233139575491367,
  0.240536124890415, 0.0906785757394191, 0.284472702855253,
  0.301798069130606, -0.39437381415882, -0.510589973915199,
  0.815824110549077, 0.625739784685856, 0.145219495267664,
  0.0242960652739215, -0.177597040482814, 0.0309770924205433,
  -0.46225387985027, 0.127137546096095, 0.843080466817099,
  -0.0791973917786961, 0.681566705090969, 0.693282340655807,
  -0.0342276027197955, 0.142664669382977, 0.291222487649876,
  0.560938624743593, 0.423459524134432, 0.426280032036736,
  -0.735287985008972, 1.71047332086016, -1.54550787826394,
  0.142107582400246, -0.0778484181959115, -0.106608605669041,
  0.228232663674004, -0.138865384396477, 0.319458332674039,
  0.39580302988468, -0.299563521963809, 0.455553755708455,
  -0.140542649537691, 0.291799017972747, -0.127168985659593,
  -0.498504982562862, 0.531536785885102, 0.290780428109606,
  -0.926489767416198, 1.85981038438844, 0.627539456954857,
  -0.144568552349074, 0.165167922159542, -0.113733890111684,
  -1.4337130342366, 0.200098127921642, -0.203443951502961,
  0.13057232570401, 0.177300240803046, -0.079411297891389,
  -0.0358905625588208, 0.201180640856806, -0.153165687335145,
  0.9106949914044, 0.816182877092826, -0.345330489392045,
  0.660106101531777, 0.176832218334768, 0.326762069579135,
  -0.0492372813916094, 0.112918516525408, 0.220559655663305,
  -0.150552081002479, -0.0951718500975187, 0.553495042975769,
  0.947834710993144, -0.147674044162065, 0.733858803201193,
  -0.148097811665198, 0.0762575014902344, -0.457676741049319,
  -0.202333841833426, -0.893166160250022, -0.35092234565728,
  -0.167436155208072, -1.42643033579979, -0.320522503709694,
  0.0775310653572296, 0.224557102515786, 0.158173902793332,
  -0.218524757977496, 0.175124436962018, -0.116902260407649,
  -0.319540102925718, 0.20390909641228, -0.0478167726178325,
  0.163439472044364, -0.127702224603302, -0.174594410486922,
  0.102384410378039, -0.108556498483469, -0.193778786719378,
  0.218276611948825, 0.203465180622056, -0.194803210407764,
  0.171965346190744, 0.10103436896372, -0.0210635707390134,
  0.108384181394318, 0.527701287428942, -0.062349650388096,
  -0.826726545379917, -0.346298175841075, -1.48170817824667,
  0.0414535677416919, 0.00314354008614713, -0.345178048887957,
  -0.0307915880691106, -0.643718519179544, -0.0167090796301592,
  0.435371767455142, 0.423100378700064, -0.180503463345557,
  -0.253580043855046, -0.0473898601193027, -0.321305125049666,
  -0.234222633527051, -0.570972404359655, -0.348029953005529,
  0.217841631949929, 0.975844283631728, 0.906115686391732,
  0.381099483209079, -0.147961491544131, 0.238792309738896,
  0.159118544603382, 0.598823600883993, -0.143778666521256,
  0.387538888412975, -0.117834039310643, 0.981251808238531,
  0.14330960456721, -0.213046683351642, 0.1304930824789,
  0.457589761249406, 0.0146366780758045, -0.278773118215352,
  -0.270455805742164, -0.314230650366444, 0.958237105613589,
  0.102652788697308, 0.173304901460874, -0.195044936480953,
  0.0995156560987546, -0.155907357094385, -0.69166578533968,
  -0.0588376740197107, 0.227911452161307, -0.0538330219795878,
  0.0988251589341292, -0.0908645343087043, -0.294204838643021,
  -0.375987027743236, -0.159713844564889, 0.595354402922644,
  1.61006817107812, 0.120839327387443, 0.328697849776409,
  -0.0926025969290744, -0.111129945825893, 0.252419344777164,
  -0.262704230107182, 0.192974554616405, -0.382111753523452,
  -0.13514611076548, -0.27116068724166, 0.755198357993374,
  0.600632814854038, -0.365215081370871, -0.0487184193109994,
  0.775824780714394, 0.444132297376494, 0.854057517067136,
  0.783255088235028, -0.0804915883689352, 0.188686218297478,
  -0.0359142397880412, 0.0581216824277116, 0.287915803374178,
  0.138276180063949, 0.00272351130450619, 0.201594875904634,
  0.32017657731338, -0.336465160374109, -0.832092454944557,
  -0.204096951287237, 0.122717730263246, -0.00768156792007888,
  0.0794996079935841, 0.561596798960511, -0.332309846458551,
  -0.28512144629851, 0.832566564117782, 0.711229503103711,
  -0.0323242423239256, 0.019715351836623, -0.206379423266918,
  0.812621190612796, 0.788847029756517, -0.150312896212218,
  0.297901938940021, 0.722044274547911, 0.693956048653977,
  0.255265071049222, 0.0688571537347121, 0.225599110881275,
  -0.337780255241389, 0.365571792691207, 0.0317071587399223,
  0.241503441059491, 0.604283552224417, 0.316712142568356,
  -0.0876906661376483, -0.0875393425685733, -0.15165803734216,
  -0.0249471572411821, -0.00267706841177951, -0.414610910278561,
  -0.0425020209739507, -0.225282553933174, 0.0337450884057649,
  -0.144318847853247, 0.0963686976583308, 0.0728224401242479,
  -0.680978804355645, 0.29196500266826, 0.506427190115098,
  0.623400908385118, -0.00481807032531437, 0.561441274085412,
  0.0665310314222628, 0.228032627271971, 0.140516147825369,
  0.85387043219528, -0.665180803942944, -0.177245330914215,
  0.404689756186127, -0.118529804599791, 0.675607161875942,
  -0.232938962520253, 0.0283620168640032, 0.185866641047844,
  -0.650736593176999, -0.241621054522846, 1.08536686592732,
  -0.26260662392989, 0.0096557572714473, 0.241666989198709,
  -0.0900075131202738, 0.118030496057578, 0.0355199926074972,
  -0.77388758684124, 0.193153757995134, -0.528362314845239,
  -0.0309886916380043, 0.672480941377076, 0.0795281497723401,
  -0.0621062309541831, 0.69848769361317, 0.00909605958141125,
  0.445652628605708, 1.42821782258981, 1.07084276099635,
  0.703811046622545, -0.00764000744907406, 0.755299600755916,
  0.080042154150812, 0.324449077347298, -0.196339320889035,
  0.39708595921804, 0.503545697941748, 0.42117062954472,
  -0.612464894293067, 0.0642309774567622, 0.00310762387992573,
  -0.32583077031104, -0.144888095154522, 0.310046508478182,
  -0.305226533695386, -1.09981421050398, 1.31273949160975,
  0.622407770146858, 1.04456296130784, 0.365428457354941,
  0.014351930595564, -0.145822110625208, 0.0758469320127121,
  -0.651782926046207, -0.943461885507269, -1.09991947852481,
  -0.144272372318107, -1.38560912086229, -0.247818112330218,
  0.13516598487604, -0.0455440497259268, 0.0967245083066104,
  0.876658733313678, -0.914295365824379, -0.741734808571426,
  -0.447164999965743, -0.235153812210097, 0.541703161724548,
  -0.210108673904278, 0.198098375394395, -0.378999270518783,
  0.625315829250857, -1.25293634686545, 0.163337252337491,
  -0.742911770991267, 0.464443904727239, 0.440023888107528,
  -0.0248023360695869, 0.355900727949995, -0.123659963816699,
  0.428606656334645, -0.965078265853601, 0.0775159356711056,
  0.229462543805428, -0.0692507389271134, 0.241837728052645,
  0.0212942478626313, -0.0353762783035835, 0.28084148501635,
  0.142018098850547, 0.943753402027375, 0.173472639016597,
  0.618266765853931, 1.23694675118046, 0.255607025261886,
  0.0106975536635057, -0.293247071986466, 0.0299335470124737,
  1.67509210236066, 0.208551860048046, 0.201623952392309,
  -0.499413823587376, 0.00672729244361203, -0.979305269380394,
  -0.135398987982775, 0.0540736190370174, -0.218036247457538,
  0.179231152012346, 0.150619367684075, -0.966469192218274,
  -0.204464323877621, 0.785793818673188, -0.161947873700527,
  0.00522034982952793, 0.230387410306072, -0.228693953014438,
  0.382744502760646, -0.641990913322134, -0.458474492034989,
  -1.43791324186328, 1.4834531416026, 0.430822063354803,
  -0.103421848537645, -0.272302084788332, -0.165081363234752,
  0.48639565636749, 1.02822488647646, 0.630701138946614,
  -0.135938781731159, -0.245834823536479, -0.26982136753134,
  -0.0567518592260814, 0.0812567813113021, -0.0776026995731899,
  0.373332918178697, -0.719233084319006, -0.567669317930365,
  -0.542685213291881, 0.0109900966688451, -0.509514058237901,
  -0.00845241044242665, -0.193124432595316, -0.0206237639335843,
  -0.0226993667931639, 0.574295058162605, 0.452633412808965,
  -0.268590819044939, -0.90570949614228, -0.948393917247048,
  -0.193843228148696, -0.0896755692505604, -0.0423849939631468,
  0.138420494794712, -1.23416238488355, -0.32338820897585,
  -0.947074250330442, -0.13888044411164, 0.926069625373203,
  -0.624156526989596, 0.225127186729957, 0.122916460090344,
  -0.927588539699678, -0.60151714153785, -0.103460943639335,
  0.346916721976186, 0.336574390113244, 0.220581933432842,
  0.14525151230141, -0.114546937729996, 0.0187350589842819,
  0.328170043719226, -0.110319390645798, 0.298660238436016,
  0.406019183655304, 0.523097952892223, -0.319521241036976,
  -0.086419201535037, 0.223442867862684, -0.263671677235745,
  0.651130143270037, -0.542617798736669, -0.301296049945797,
  -0.289907758000346, 0.591924580164066, 0.83668093966777,
  0.371411141988112, -0.0206260276174877, -0.0159925990372565,
  0.85349654180487, 0.34634772077242, 0.357735036394028,
  1.84210948833196, -0.746696615111111, -0.70612171628896,
  0.0559321820927432, 0.316900021325738, 0.179697507792565,
  -0.128776277783351, 0.183712738563994, 0.681782087072308,
  0.205895990978263, 0.362414797185061, -0.156016469990143,
  -0.0646496141610429, 0.0938685569591526, 0.199898070266939,
  -0.0915650569103626, 0.368784201262077, -0.024611766183373,
  -0.949399954360356, 0.263233538693823, 0.140380142197338,
  0.132347915568627, -0.0454118209718935, 0.00508474221172343,
  0.0627447080042013, 0.679491879446776, -0.891446475205536,
  -1.20061690989169, -0.51572513476383, -0.796391509711102,
  -0.117591929679698, -0.0484930117179008, -0.13682837589241,
  -0.561696103465118, 0.15343769445092, -0.550345455318976,
  0.975961026861437, 0.20460294342425, -0.0343573776380034,
  0.0592368296020746, -0.0290657120583858, 0.194906685082129,
  -0.0156053492643795, -0.339397208396664, 0.286474086171109,
  0.0473368189117214, -0.615726757148065, 0.263785815271404,
  -0.308425408313091, -0.206241690529445, -0.131148927736987,
  -0.793171535434894, -0.170017384880783, -0.386778055291622,
  0.0864985716780867, -0.210503441506617, -1.72060922465424,
  -0.111000789141957, -0.109531490461006, -0.0747866263309283,
  0.41028045148949, -0.302095831749318, 0.562985642608642,
  -0.0880551427451137, -0.613872912425367, 0.150849198834356,
  0.104151676133479, 0.253052649200945, 0.270885891657583,
  -0.150023756764995, 0.119156749493444, 1.08000220714377,
  -0.0663384402062792, 0.660590202955121, -0.17529742329198,
  -0.211275717198591, 0.0821001293107169, -0.111764111423388,
  0.0882893221891513, 0.685591279206194, 1.02519366055723,
  -0.404373575819945, -0.485932044376703, 0.495150207915739,
  0.148082148242658, 0.00522032809779286, 0.124624745775447,
  0.654273452208391, -0.490177051368823, -0.582884250295815,
  -0.171938213396284, 0.462397416835474, 0.703251369331781,
  0.124841921168735, -0.199453517390698, 0.284162863357855,
  -0.409501557677031, 0.613533824213489, 0.553019607774526,
  -0.532049074852448, 0.50585901779718, 0.621619323391547,
  -0.0083120499963383, -0.143589174693959, -0.659908217070859,
  -0.0308736612361135, -1.08482455660442, -0.865818715792204,
  0.593357141088174, 0.202987914611493, 0.250772916984866,
  -0.16752894615054, -0.0458193469027414, 0.248545210027405,
  -0.81009297503875, -0.646510472100324, 0.498021742687783,
  -0.291184069710436, -0.133846094084348, 0.245361590753466,
  -0.10377376370505, 0.012223542907096, -0.219534554149802,
  -0.559411773044548, 0.719599270679047, 0.618356921014511,
  -0.531728830919317, 0.717168502432137, 0.623883256250648,
  0.193282481964231, -0.0236530553567284, -0.0988990340161662,
  -0.369278252274144, 0.226794650869769, -0.329264725527866,
  0.381965819977122, -0.805960670202818, -0.347241890403971,
  0.182030415966124, 0.371356154849664, -0.0617840186074799,
  -0.711551598741642, 0.613741679684579, -0.565228278388214,
  0.161683526559538, 0.811072155227334, 0.740458356124983,
  -0.0849232371526338, 0.00394351917044318, 0.0739413035159716,
  -0.158851986417835, -0.0197534853346228, 0.659116505921453,
  -0.421646889078054, 0.177779858876758, -0.00384880526604132,
  0.123751343015689, 0.321289298890759, 0.103205909222632,
  0.212528323837249, 0.725848638044283, -0.170774579734992,
  0.162278590026076, -0.0681379043349248, -0.227051222943505,
  -0.296808457040061, 0.103084847663071, 0.35675430821532,
  -0.15625703894275, -0.165458682359185, 0.716549360489284,
  -0.333188931943975, -0.222489785570729, 0.375995833261413,
  0.0273921816442601, -0.112808479444377, 0.240823867892474,
  0.0796085514195368, -0.593009445442836, -0.15976918391875,
  -0.307166307547372, 1.34910007284731, 1.40707826617512,
  0.0182755284733301, -0.0559321093441352, -0.332736776520207,
  -0.231383584528507, -0.0759159359631188, -0.637274791231904,
  -0.419642704419891, 0.117955817618529, 0.848665678825175,
  0.199670749536743, 0.0503583057357138, 0.178059834466183,
  0.173381611080687, 0.369893335593157, 0.0949760582024994,
  0.00746223242407355, 0.138961343816295, -0.137534156161902,
  -0.107039603670707, -0.325660736700393, 0.348785781631452,
  -0.436598363015319, -0.267605508228586, 0.0176221803437846,
  -0.833953979435372, -0.218533670395751, -0.125745296925531,
  -0.150628378176896, 0.0239635844498329, -0.186021519768128,
  0.880556402339158, 0.02967633742524, 0.210696335300289,
  -0.519022314679514, 0.0244705835371479, -0.33474430658339,
  0.34910234945697, 0.0700645895721552, -0.0815605020275073,
  -0.819861362718893, 0.288233029130225, -0.570755504391363,
  0.0256437080365621, -0.202220641429346, 0.569362022791284,
  0.0771574696568856, 0.0119046901234239, 0.192188901694832,
  0.342767031363346, 0.534286004527483, 0.0927845559175849,
  -0.141711046363115, 0.0906307610000219, 1.72263934150896,
  0.33897595114777, 0.183724031037498, -0.173391299889284,
  -0.444539860667391, -0.46421478409427, -0.279851581979143,
  1.13192137967305, 0.0844159400171307, 0.0208500565725315,
  0.200252729334734, -0.041236480410892, -0.36035668107947,
  -0.341251156770587, -0.735094479538871, 0.697340698050973,
  -0.523348081129594, 0.530253603598355, 0.331082339659708,
  0.396390520154871, 0.0523578605466507, 0.093310100956746,
  0.497990814608673, 0.466734703004338, 0.398258725480165,
  -0.136786993206631, 0.0263784775631447, 0.0179932159145792,
  0.278756770980599, 0.507276013502298, 0.0993588281580993,
  0.103766727708077, -0.0866252568131923, 0.342929919023131,
  -0.0327673976991207, 0.403474571493486, 0.213569520296113,
  0.103783509213663, -0.0326848318592444, -0.299437599191645,
  0.454379706137631, 0.266913698071952, -0.0420446678812652,
  0.439393038603341, 0.689142049666112, 0.465989913841997,
  -0.199425292803952, -0.127239037279515, -0.120787190022777,
  -0.55939338423891, 0.181091725802886, 0.0593311195342582,
  0.0248771333441378, 0.347098182150005, 0.18872414351791,
  -0.114058296027475, -0.0471023052534609, -0.133176970064667,
  0.028966616295551, -0.57125382586766, -0.286223173032883,
  -0.201994214668901, 0.2844146225583, -0.489782511277327,
  0.34427278113805, 0.0355509513544894, -0.0507693949326077,
  -0.487940244601789, 0.373226115133015, 0.44207092366563,
  0.475743393889783, -0.960853124314266, 0.149498675472586,
  -0.210888013369974, -0.00568025875042607, -0.108532709261702,
  -0.0920601951938476, 0.313092387940593, 0.330531192952587,
  -0.227634026649927, 0.326368367556122, 0.509137050963049,
  -0.160428513798104, -0.0931118364052898, -0.496348853019583,
  -0.236740471290717, -0.413681200671692, 0.148439367544951,
  -0.475265814237248, -0.160158799760574, 0.255567923559841,
  -0.00425439579171922, -0.0060831710116169, -0.180300744257033,
  -0.238073972034609, 0.250858810623031, -0.342494734158729,
  -0.230164391817657, -0.205981256944017, 0.0623482435638477,
  -0.0787358688791658, -0.0622158774551169, -0.038062130825726,
  -1.51683989517916, 0.565099695440269, -0.13380869020741,
  1.48011116237293, -0.894736602757171, -0.398408650896053,
  -0.297511592324728, 0.0810631250384055, -0.215541167343245,
  -0.0209645490682785, 0.208749338991839, -0.654900070890502,
  -0.411116863864587, 0.016490343069184, -0.031272170878401,
  0.148414653139747, 0.457024732883097, 0.0254940552427736,
  0.366974982971806, 0.648609346511687, -1.0164295270392,
  0.0603036417462688, -0.338948000070949, 0.452218787170186,
  -0.0685324566966133, -0.00427278555390571, 0.227861130457731,
  0.229960637947214, -0.371250779937132, 0.952565373204045,
  -0.684725262320722, -0.741163749544163, 1.55449707008193,
  0.00553381783177184, -0.0820349659557366, 0.0196611237434319,
  0.177968078393571, 0.0534069810684634, -0.196845968715702,
  -0.789259193303336, -0.697450900853982, -0.0113676497040861,
  0.0478923973071456, -0.0486244006117013, 0.213708680240975,
  0.0786360135896978, -0.429529544166561, -0.0919913256503892,
  0.313215017573009, 0.258056367762336, -0.215386938433833,
  -0.246440982459843, -0.228848732731333, -0.42843833179342,
  -0.749635046778478, 0.159894878644211, -0.798751983776543,
  0.167297374881099, -0.729152018465428, -0.501853842253821,
  -0.0614390794457734, 0.184038312204406, 0.304158314255825,
  0.999641119836026, 0.118337443274847, -0.354958491851263,
  -0.630102245823031, -0.718968619797239, 0.734843107237369,
  -0.0291280425088313, -0.0148625695481588, 0.199729709362113,
  -0.117141927959072, -0.0418532136130896, -0.297765985199325,
  -0.260858046289437, -0.436772068354001, -0.623911726877933,
  -0.0290273871500666, -0.164991439139313, -0.0416474807397493,
  -0.377360917933216, -0.364329379690775, 0.471779064745775,
  0.245295993871065, 0.000790901736324197, -0.302582549201134,
  -0.033488560912289, -0.01082205398747, 0.433757751858089,
  0.403516943694695, -0.024385239035102, 0.503759234293889,
  -0.239170473652269, -0.137618995725984, 0.432141632384117,
  -0.178653596015348, 0.215354952003186, -0.0876971668315233,
  -0.140384786166363, 0.650238587937106, 1.43589876924196,
  0.0755550065720484, -0.722208992234155, 0.449019661288782,
  0.0974451532656084, 0.0724116520626949, 0.0774918145998282,
  -0.100176406271905, 0.454292451354206, 2.93927160628113,
  0.512497859720759, 0.105020972897536, -0.277591914239048,
  -0.00320106174047621, -0.185850884446052, -0.119067398793401,
  -0.265194541084425, 0.0088155040707484, 0.0276238257526581,
  -0.0443022650804413, -0.304416380442708, 0.140220996458289,
  -0.215106694467328, 0.0938305984892808, -0.0658550682251919,
  0.174041617579073, -0.179034744717844, -0.0930617172388069,
  -0.491514689511457, 0.39925184227976, -0.115890060236488,
  -0.0311914856935632, -0.274108091373614, 0.0665417999023707,
  0.170577268727219, 0.251435911112419, 0.576874766532674,
  -0.799817787672753, -0.0678140776700366, -0.262793992081293,
  -0.216866173331226, 0.194381330431839, 0.00352326574557527,
  0.599510455085998, -0.146247938069849, 0.65558133355967,
  -0.551333410558004, 0.00219967294362134, -0.529752428624203,
  -0.268326031047876, 0.133493978653774, 0.315449467184642,
  -0.934247604346038, -0.444880511839053, 0.450475294041463,
  0.174713014674639, -0.128349710436567, -0.512571087098542,
  0.156240326263328, 0.0209965640749974, -0.0538925023206727,
  0.323074075748421, -0.290758475690485, 0.897822302667561,
  -0.119743497020339, 0.348306190875294, -1.73706572126931,
  -0.391479827086577, 0.0748576916941207, 0.256182328022052,
  -0.46260311753485, -0.250150986420608, 0.247063568936635,
  0.701796032382439, 0.157854975202848, 1.13396995569249,
  -0.222171094089984, -0.0702447798058389, -0.0803740390796941,
  0.15260690098994, 0.636026787778186, 0.573538790545542,
  0.743268325359123, -1.38143094625841, -0.125989558366654,
  0.00929708857968817, 0.056649535063999, -0.0469184316994726,
  0.154694195689032, 1.0270395279008, 0.6325801216503,
  -0.495659575689577, -0.333986782365811, -0.122881992403169,
  0.275836706241135, 0.133217010819018, -0.0952246107423356,
  -0.0289246530166361, 0.430354674911963, -0.36121061984984,
  0.856377238208241, 2.55012704316363, -1.01501697587268,
  -0.228676535179057, -0.0556995000115304, 0.312657764647069,
  -0.546640639301412, -0.0477323437749807, 0.560731659604002,
  0.498857950786055, 0.0542864013785236, 0.259346395762041,
  -0.0240641873511867, 0.237991744822318, -0.3702621835604,
  -0.725157027716721, 0.574139368323551, -0.948715601929188,
  -0.175144541219493, 0.126931441149682, -0.742387742614173,
  -0.0331112961851038, -0.0497446312834777, -0.187480780773291,
  1.04742089108088, 0.323031113610898, -0.078083950070857,
  -0.275473048272908, -1.51065407927752, -0.0319707812238887,
  0.0488080228764587, 0.0225654373133433, 0.213493105242117,
  0.0749042800354751, 0.732690155139686, -0.272668076739144,
  0.083907254700355, 0.180746232142296, 0.184005356122652,
  -0.0694788624028654, 0.360714393154135, -0.140010604486062,
  -0.577855959427868, -1.05316658911269, 0.378625162783863,
  0.0992505692683626, 1.20712995584528, 0.795472386139206,
  0.155002942865096, -0.0436645483114977, 0.159604405679124,
  0.730405207323038, -0.130063207184387, 0.213163448146818,
  -2.03584589374703, 0.429030443520667, -0.22488968564878,
  0.111352987174449, 0.0586724113294511, 0.0131383137931928,
  0.704167140920524, 0.608326814919178, 0.316771056320127,
  -0.231541438602641, 0.382619651924265, -0.560927874769554,
  -0.0444330198226008, -0.0448488171970673, -0.0510452806053926,
  -0.986780285578301, -0.255432981280638, 0.360519689274641,
  0.267742165880054, -1.41669602885291, 0.333745768371552,
  0.0127889753590681, -0.0488118305223111, 0.129225578357564,
  -0.464952570740713, 0.201239087140324, 0.556569549615519,
  0.444985337972258, 0.221658852097919, 0.246345937613258,
  -0.00240052405875753, -0.115603452846721, 0.173265284615086,
  0.116364536022193, -0.823261807998745, -0.397543856851156,
  0.521810991631504, 0.252721974865067, 0.147270666795509,
  0.0536468066478649, 0.0497657400589348, 0.135075738421531,
  -0.449447206657434, 0.256707068423757, -0.0244362962593969,
  -0.928867505930625, 0.427133915675173, -0.298597052911043,
  -0.350964989961794, -0.112645976699452, 0.043701619748333,
  -0.0299764340499188, -0.0414020627959261, -0.853216446522016,
  -0.643903391819232, -0.205601862885774, 0.203757516561938,
  0.124304799076518, -0.175280207555161, 0.142648141790385,
  0.341867562872869, -1.22400169484615, 0.114306706890717,
  0.411655774281061, -0.421391299694257, 0.140663536542902,
  0.120644098958458, -0.114649617182964, 0.0137619627922482,
  -0.113701623544526, -0.042022225881308, 0.661655945034287,
  0.16652013142251, -0.316820225369589, -0.0068664354730063,
  -0.215445176620382, 0.237822524388092, -0.237452515138225,
  0.142503080215899, -0.00672660404011829, -0.265241132653573,
  -0.553205070731243, 0.360316928077862, -0.262232234193219,
  -0.0736521425502438, -0.00966345179435526, 0.425679493842241,
  -0.694798817113304, 0.38160351533558, -0.438277840049496,
  -0.236314921550715, 0.106288236865935, 0.569858570922863,
  -0.263571205174036, -0.080931667238503, -0.0801891611752857,
  -0.442591823468131, -0.00888178654582176, 0.738631425909801,
  0.193752169390325, -0.00570804274896692, -0.888666781203197,
  -0.0964079942170373, -0.0363231640735063, -0.0967309728053151,
  -0.257868234579765, 0.406813558508108, -0.164380405183465,
  1.62238677659659, -0.406892138250348, -0.55860525899076,
  -0.162202450526753, 0.161907139313263, 0.211474559995644,
  0.498488563211235, -0.0315450595752817, 0.720263623157887,
  -0.570556871933631, 0.572845581358442, -0.497157402106709,
  -0.196842628197595, -0.00445775018829642, -0.0202605813332106,
  -0.689151119359771, 0.0292260493512894, -0.699471575284576,
  -0.388175359532593, -0.112943431920937, -0.506290873967907,
  0.300885006890303, -0.169418663964531, -0.355081581618676,
  0.425965166877602, 0.218827449687787, 0.143183429945076,
  -0.00447409487670639, 0.221525368314236, -0.487141490732376,
  -0.145043867694368, 0.134028917447619, -0.188649457895406,
  -0.104054987415324, -0.383928928405777, -1.26380646923586,
  -0.997938841220552, 0.0984305272781033, -0.137484991426065,
  -0.280373861040143, -0.0633281326806848, -0.244924786622438,
  0.478988852560054, 0.0933911641363267, -0.0420505282119601,
  -0.903282184239975, -0.152674514147632, -0.0912414889696986,
  -0.0489492942460416, 0.077279065657999, 0.190921573234737,
  0.732433254969671, -0.145100689678511, -0.261962483502384,
  -0.201205723252545, 0.772466048104895, -0.0576750001273185,
  0.105717447541137, -0.0644141557376277, 0.195531923511269,
  -0.236237280192183, 0.183519328642373, 0.516693986322662,
  0.172824372468813, 0.445610216226844, -0.0283640395143467,
  0.103562634527339, 0.0275811373988801, 0.173341407392339,
  0.352651998036169, -0.38675305790714, 0.691343865115836,
  -0.307090906434621, 0.39631294430029, -0.689303384808256,
  0.360695493684135, 0.248632730158507, -0.104915170091253,
  0.625645557013808, 0.678283569268304, 0.077432013393206,
  0.124151317248668, 0.431660661147114, -0.252633685459253,
  -0.125021539638766, -0.108729634091495, -0.261441648241297,
  -0.0644289852941951, -0.125185024850229, -0.031736712967284,
  -0.249465818607739, -0.375514995152085, -0.407246396621019,
  0.181896469178092, 0.273979422516172, -0.0206378305163399,
  -0.0389316999219737, -0.0637720151178658, -0.164966852572141,
  -1.77602861704071, 0.1763553009178, 0.532072791720956,
  0.246903001281339, 0.36465104540401, -0.0025179098576035,
  0.516357859530633, 0.782530642481467, 0.0425522042569938,
  0.403735210863558, 0.0610777755069541, -0.391444575334838,
  0.391940620299381, 0.163323307698376, 0.0966612835039608,
  0.274409782465267, 0.667308996326492, -0.421853200700828,
  0.731589072520769, -0.311043919097409, 1.26447884492489,
  0.0540285495355146, -0.337986987237402, -0.0476468613577362,
  0.135000116223806, 0.081074773754268, -1.23850901945763,
  -0.0957268461524551, -0.573890975915769, 0.47766321990558,
  0.247609195842968, 0.365233967401045, 0.0284874370928324,
  0.44389884153669, 0.256212139764447, 0.314201558754074,
  0.273821392954655, 0.330504187587566, -0.50142582490859,
  0.0631278500313912, 0.261549148345207, -0.262442144553293,
  0.100955685146421, 0.307318340955345, -0.268064521949179,
  1.39269299284913, -0.22736104362915, -1.28370377191742,
  -0.0523828767156289, 0.0737652267047345, -0.127141000065002,
  0.202835126353965, 0.258813715682469, -0.991692280772975,
  -0.357612960759547, 0.76063357406756, 0.267124018613575,
  -0.22997509824064, -0.0882207026105804, 0.171161741186243,
  -0.926150310082232, 0.141046674742609, -0.370455605989748,
  0.452068351446795, -0.0459756344432541, -0.20556622991685,
  0.439702340800211, -0.0236831047923426, 0.152282606232663,
  0.0778377678463557, -0.0015726360782348, 0.18721065580446,
  1.31749303946907, -0.354255029370178, 0.606297170109208,
  0.0930185002035006, -0.0091010045087871, -0.252381565723241,
  -1.30048771299459, 0.203961225277416, 1.25140905969975,
  0.380537154631786, 0.178097146593095, -0.230194215485394,
  -0.0342261445096819, -0.13748693038054, -0.190604941892933,
  0.0481947807369813, -0.554628456289172, -0.322397838829828,
  -0.106630002053822, 0.257917459503942, 0.244525752780525,
  -0.397046337040489, -0.371897961461668, -0.118519456496114,
  0.610746077923158, 0.678206292875506, -0.325262233932989,
  0.360592819800117, -0.158538713291923, -0.798142164870223,
  -0.091730683786644, -0.405907909930656, 0.00479772742808424,
  -0.280431768518809, -0.234462508875751, -0.694032004634492,
  -0.101585607520777, -0.47265847067529, -0.505271963755592,
  0.250116607216977, 0.0533465879856909, 0.200269478490738,
  0.259080114819945, -0.167702804150136, 0.250124263748992,
  0.412848338606004, 2.0620782160472, -0.51074017978861,
  -0.138644350654875, 0.248767948458293, 0.144267423791248,
  0.162332800410811, 1.20773066815931, -0.235624348803778,
  -0.941258095244087, 0.314139782355015, 0.0419344353309877,
  0.0838531489951432, 0.0483579333609977, -0.160555577050215,
  -0.134019200340367, -0.127349763451216, 0.158477589830575,
  0.135810502157346, 0.103102850031322, -0.283706016805285,
  -0.0838022460701274, 0.163981917207542, -0.117649454489763,
  -0.683542563799665, -0.167574145234648, -0.514328944705106,
  -0.489533927633226, 0.22012269158322, -0.192759896468954,
  -0.281633318310327, 0.173527414872856, -0.182016704470978,
  -0.779357905786057, -0.61307247579243, 0.19678542311804,
  0.133563245164832, -0.0635320618674299, 0.566413669587476,
  -0.149380005594837, 0.109797135278819, -0.296791441317115,
  -0.187871012983562, -0.108829620017441, -1.40481892212223,
  0.636849866591668, 0.2916678754114, 0.124460686668985,
  0.11965160137532, -0.149611714687338, -0.0950602862058703,
  -0.887768960755046, 0.0623277201354063, -0.185558296943994,
  0.310247545718564, -1.06561213636107, -0.289392690475172,
  0.0360354435945751, 0.247163031883588, -0.0561534127581552,
  0.222435785083896, -0.489153923359718, -0.313718674980747,
  -0.150492728005033, 0.048668079788623, -0.70193717773227,
  -0.237906296956886, 0.616351606347504, -0.220630347477759,
  -0.0369413636487656, 0.0054464789336168, -0.370300224057228,
  -0.294407958349816, 0.853344025428091, 0.298975162988515,
  0.193060127476092, 0.0539087171978662, 0.278859029150743,
  0.431836056927883, 0.0374442277909009, 0.74331806162594,
  0.00118809612351761, 0.703075484951405, 0.0909879468587823,
  -0.190651277945373, 0.227069370865411, -0.0283576060912485,
  0.126110818376102, 0.521127057957074, -0.00434065992503374,
  -0.574095535399818, -0.0558692519137906, -0.0069833494884968,
  0.169784789960659, -0.0845248822055606, -0.179387594497375,
  -0.0210022055003454, -0.663192941184043, -0.297530774446275,
  -1.22438617730387, 0.0137298661335351, 1.09973996829887,
  0.342730680334453, -0.0489971898969732, -0.0243759336993502,
  0.245106560159208, 1.12981885898029, -0.416029861244966,
  0.129385692871178, 0.494851689261189, 0.0662722175526738,
  0.012159323639185, 0.197679651856898, 0.193117192557799,
  -1.61994065263172, -0.253151720412887, 0.523197549825265,
  0.233348251925983, 1.55830114777818, 0.606947510566063,
  -0.111964112305883, -0.0122983504615814, 0.229256832442896,
  -0.16179987287025, 0.658132727186343, 0.110799614523757,
  0.786587178161095, 0.278110094607832, 1.03530484479915,
  -0.091335198652641, -0.153298580922944, -0.101810286814085,
  0.576865440346375, -0.0491304721762248, -0.96413664933246,
  -0.56631176913739, 0.813829320887093, 0.426906161658066,
  -0.0236195467151026, 0.104326106896414, -0.181785774472695,
  -0.471650060335524, 0.498294057063666, -0.204533943913129,
  -0.117598123696615, 0.188900408397744, -0.20467829888899,
  -0.0776631039582119, -0.120425715464579, 0.190839863259695,
  -1.08285834135139, 1.16824233633569, -0.0912057240555417,
  -1.2037268153347, -1.25535374682381, -1.57247653609766,
  0.0116971381905984, -0.180971723134545, 0.0669783963499721,
  0.0411252227616865, 0.548963502546253, 0.107628794662712,
  0.0845618241171724, 1.01088666853417, 0.172388513337045,
  0.240539780505176, -0.253946092950934, 0.151076444329349,
  0.131465968927214, -0.0445410945041984, 0.480965141071335,
  0.0905544369684435, -0.0780205271517066, 0.242554451927321,
  0.161065375540197, -0.249772261325802, 0.0157407948899034,
  1.40592916178787, -0.90922761159074, -0.431284752447579,
  -1.1171656610385, 0.748509256365979, 1.34466902936786,
  -0.159076236145202, 0.00701192120529189, -0.213103506433714,
  0.271718083212393, 0.541328266097602, 0.785262705008133,
  -0.443461640825118, 0.206670903187951, -1.74460030538639,
  -0.00550258359297997, -0.107719929221804, 0.140393489637898,
  -0.157113811420294, -0.899226460813617, -0.0707246763469329,
  -1.43169854327846, -0.50910626592426, 0.92651719339195,
  -0.316092061741583, 0.357919004880373, -0.368098564223658,
  0.0273610376927993, 0.125757940603254, -0.453808130708714,
  -0.0241913174840884, 0.340095635628897, -0.164359334944053,
  -0.348573358487622, -0.120596091867513, 0.000822558119219611,
  -0.545288309354471, -0.339925518391997, 0.200160381474942,
  -0.485951945583391, -0.228937956127207, 0.0237679819617817,
  -0.233155891256424, 0.0196992082381142, -0.196115448766804,
  -0.378543905747249, 0.457333506916582, 0.497861410906144,
  -0.838783353169706, -0.128395219228077, -0.876952101093765,
  -0.227227375242782, 0.180630836117297, 0.160548727384201,
  0.341432493311113, 0.301100869864026, -0.443571851611703,
  0.478923160280909, -0.298816854303025, 0.304881535139445,
  0.361619464458558, -0.349163554915836, 0.292381989968029,
  0.495918781961472, 0.265721302589771, -0.00601247718885021,
  -0.615452460425214, -0.823816153695965, 0.263295180821494,
  -0.138106000870536, 0.386769912373044, 0.431275686408587,
  -0.0988795141938559, -0.507255374162504, 0.341701184371008,
  -0.210229779222398, 1.10951712991139, -0.585168957533435,
  -0.0381102157931578, -0.0123352308125939, -0.0520807237010727,
  0.0261763704091006, -0.273937704611102, -0.146509032921151,
  -0.261537697944722, 0.0661483522523546, -0.161571182419714,
  -0.0778960601160578, 0.0261348091692385, -0.00365245449781034,
  -0.271806913167192, 0.606263422137214, 0.23636887097391,
  0.514729356105251, 0.193746685916056, -0.472367788544208,
  -0.132652293617019, -0.0908859455827509, -0.0205643569098803,
  0.172938704910771, -0.235395884761167, -0.565983798891127,
  0.368158950796784, 0.0959797061044819, 0.544095741858899,
  0.127780348191262, 0.210192870633217, 0.0393160579048031,
  -0.189466370053163, 0.313289387164436, 1.0930037002499,
  -0.684183860816904, -0.194739366200513, -0.21752959426472,
  -0.335121810013682, 0.00255539931811961, -0.0188558901143641,
  -0.907449596396961, 0.0211587041369217, -0.844030577674934,
  -0.318338905969731, 0.0349483423076801, -0.957782102035886,
  -0.197084049734704, 0.177966203791563, 0.204595288315058,
  -0.45269980088118, 0.324439015923994, 0.110776084437151,
  -1.21800632807678, -0.159873146823164, -1.30525733990079,
  0.164871067694949, -0.260496620439978, -0.0229722361996171,
  0.291913914971911, -0.295745641661761, 0.488916964625077,
  0.614650522328352, -0.347279036007221, -0.534816896025399,
  -0.0573563232140893, 0.0594710568073151, -0.161988708870835,
  1.37397114539271, 0.0696080790519357, 0.445348787113911,
  0.174630828957801, -0.204345686863212, 0.138196145766305,
  0.292648213989504, 0.0433122550282425, 0.165139303381796,
  0.470869981094537, -0.044253937413556, 0.263131381739285,
  0.257637803764154, -0.114787105113823, -0.05073200146909,
  -0.0235430285842246, 0.00947345794412559, -0.0358566094075821,
  0.125437994574617, -0.489656083346794, 0.0196062569116935,
  0.0860558129838795, 0.314577045958303, 0.0782283277458751,
  -0.116155314868295, 0.0513258240297947, 0.0329011956078246,
  -0.355463392954161, -0.297038361151801, 0.990951116316916,
  -0.00410519670838597, 0.342663507364271, -0.455932642595154,
  0.195920566576992, 0.118699398170516, 0.140577574992761,
  0.858740851067906, -1.02654105581635, -0.128108829947791,
  -0.0538662637537111, 0.501133030095138, -0.330551120405154,
  0.33735119171464, -0.0181875601910613, -0.0713484784167977,
  0.361838092803536, 0.573037924079805, 0.706108633705941,
  0.0200265740714284, -0.832667657098054, 0.0940472818927749,
  0.183657564083533, 0.193116055406143, 0.109383913867794,
  0.178407120949412, 0.488197178151767, -0.984668087527909,
  0.503077991937455, 1.42422391978611, -0.0387293532458144,
  0.101605992746624, -0.225410772524843, 0.0641722379498347,
  0.162195345674638, -1.17120383969338, -0.226369507684841,
  0.0873694144131568, -0.368657419527722, 0.737151499834027,
  0.200656005626368, -0.0217992306047795, 0.093519461987911,
  -0.52063206473503, -0.252488156050734, 0.155039577676481,
  0.392619187966404, -0.621467029933765, 0.197351908841109,
  0.311401582747202, 0.0504021591703322, -0.0111951289010216,
  0.383681875940999, -0.427364245909387, -0.628148759783792,
  0.727229520404087, -0.429401284483776, -0.400837522288428,
  0.178224765385133, 0.26176792987567, -0.234240773169858,
  0.326520953549871, 0.513094156351235, 0.152513263429083,
  -0.0672490350962591, -0.100935059573958, -0.812887006194645,
  -0.0874000636901296, 0.153712817499107, -0.0925248053895806,
  -0.420889402467222, 0.522024899651425, 0.115630992087953,
  -0.327967413653144, -0.108876469488244, -0.508451316553008,
  -0.0780652302585303, 0.0368503762587757, -0.0777061935133195,
  -0.730835770823087, -0.264914059578325, 0.568455328913849,
  -0.351607701440096, 0.0138100218482089, -0.828288018304033,
  0.370185450787593, 0.140064603877815, 0.00416703616859052,
  -0.213121788102828, -0.842968975064036, 0.254122712875019,
  0.471268959512032, -0.313554645457249, 0.011420481201008,
  -0.105934507330546, 0.0944883572242796, -0.179478962719861,
  0.586127972712576, 0.254067648839578, -0.467961880366929,
  -0.545901526988865, 0.0591388014864951, 0.000825301730538353,
  -0.100984008544249, -0.1145441145677, -0.175189563730734,
  0.516472735980592, -0.540781036138425, 0.450851949773603,
  0.673542933748953, -0.633245264368378, 0.627534020845443,
  -0.0345494706455405, 0.168749450835392, 0.163007274802182,
  0.444573266325152, 0.164676491197044, 0.364783607277609,
  -0.12814781363322, 0.496391412489836, -0.0122601674053209,
  0.0678793790738657, 0.246148338321637, 0.0969906953763893,
  0.39305033171652, 0.196648921035527, -0.0949393890378665,
  -0.118549545027991, 0.583725955546347, 0.312713698305491,
  -0.30207423695946, 0.284089896133371, -0.265768219813282,
  -0.0889344322566052, -0.490836657077076, 0.0107014997866862,
  -0.489532076222466, -0.379371800217662, -0.00616539410428772,
  -0.110706451738315, 0.342024235025618, 0.31321238303647,
  -0.393543971357517, 0.152986396803774, 0.0918500653578741,
  -1.1215239672282, -0.256714396601485, -0.451356783241291,
  -0.207241259455609, -0.138900823327313, 0.055080591039939,
  -0.871962459807763, -0.255220464433486, 0.352463986108385,
  0.686577015694408, 0.583709102953054, -1.28270099246922,
  0.0349979945631533, 0.0261378247950657, -0.0793107488231567,
  0.118342991580547, -0.288306532448695, 0.0217146114023009,
  0.0581205921779981, 0.409169276038297, 0.031053957374707,
  0.0556821905521972, -0.131950606233474, 0.0613480777829234,
  -0.11788410005852, -0.750980657884764, 0.356560650566279,
  -0.423672644197195, -1.54008223257543, 0.0241653607188361,
  0.069535892389997, 0.161400659852138, -0.0622137994742756,
  0.20581567215137, 0.451172493411646, -0.126826141948509,
  0.0907685173932831, 0.237747611829293, -0.052555262172026,
  0.195280563038801, 0.0832575123720261, 0.108972005602878,
  0.756456217705046, -0.11203873618607, -0.711448620697744,
  0.517352022695505, -0.0214055596522494, 0.970611764233388,
  -0.166621016891564, -0.370877759615702, -0.0868732103068838,
  0.245261643213849, 0.25157052711599, 0.920625350272291,
  -0.74810829630376, 0.233150795168892, -0.970348889567601,
  -0.0404819932848993, -0.0560229328466008, -0.474893853515984,
  0.147299379849758, -0.108379662745597, 0.212042831701834,
  -0.0901514018008363, 0.129815247508705, -0.63599477375756,
  0.372739192726484, -0.319208130527523, 0.101256247575892,
  0.584151519849121, -0.230048261089819, -0.417921344915534,
  -0.580790201901915, -0.175069862818655, 0.235483838252823,
  -0.151497490649394, 0.311107929837722, -0.136399511180069,
  -0.98239032389523, 0.0789889897228024, 0.304888044536948,
  0.550099480003616, -0.0653164852688117, 0.309791120766986,
  -0.100828553656654, 0.273496073126847, 0.444587897270023,
  1.81725230315745, 0.930868553255944, 1.35372898560592,
  -1.88518430478629, 1.86665584250238, 0.774192564996683,
  0.406354081282824, -0.225073535964235, -0.24650007790995,
  0.333036187811828, -0.0300772001716753, -0.431335044638795,
  0.932856444170709, -0.044503648788152, -0.718918443291468,
  -0.354745302286443, -0.198356936933537, 0.103068455559568,
  0.674706364594595, -0.27462764871152, 1.26907606403889,
  -0.790758698240524, -0.134491227891068, -0.519674991691676,
  0.258142136010463, -0.0986889550318483, 0.0136030179803039,
  0.496886251270244, 0.051933734536953, -0.225427428913249,
  1.66846154753674, 0.792003568788472, -1.39122054028409,
  0.166178360257014, 0.0761149183915021, -0.136131436859458,
  0.851727477149827, 0.0486153943161359, -0.391836776096203,
  -0.353960996184687, -0.0660814261933852, -0.24084313763431,
  0.227802768417731, -0.0833382933975028, 0.0195073550889018,
  0.747458739725171, 0.143222950988435, -0.147408747380624,
  0.247272107070385, -0.366387193862642, -0.0203920543724831,
  0.142188255785923, 0.225423130391397, 0.282452702413783,
  -0.179600560187391, -0.0589133967425148, 0.731945944973974,
  -0.528473963081315, 0.293423080798967, 0.112031244458112,
  0.286256544527864, 0.00155039379537749, -0.0204273804241138,
  0.329316943782639, 0.524077112671115, 0.424661839635356,
  0.0867257254508875, -0.418812173953697, 0.296256931798115,
  -0.103002681814162, -0.0162821094211891, 0.177996296668329,
  0.129529459277622, 0.580178177964641, 0.194430349110697,
  -0.177185497935686, 0.763182280738993, 0.192148314199122,
  -0.0857185236004172, -0.169611810081768, 0.104391700480207,
  -0.805799887432619, 1.09978160479109, -0.230626753380278,
  -0.356950087781442, 0.604639067242542, -0.0887438010638706,
  0.223601941154923, -0.120130894818061, -0.306076458911966,
  -0.65563562333733, 0.416709756459138, 0.296873392387245,
  1.25899996441967, 0.372882280486284, -0.272119483770205,
  -0.187163237095049, 0.151109117150749, -0.153690451246245,
  -0.258817794978179, -0.975565204643685, 0.613927598304918,
  0.183301878049747, -0.424197652357838, -1.09530150676404,
  0.138135252197055, 0.123973295917614, -0.38426979944669,
  0.141473795472355, 0.151118579543888, -0.387510041278978,
  -1.22541816716715, 1.23958342440114, -0.530487728093436,
  -0.276568964096453, -0.00752035458277957, -0.000370960360948977,
  -0.934667023753697, -0.738308704290146, 0.634240324937653,
  -0.643423837977081, 0.400851457428767, -0.227262488090255,
  0.0206048463723109, 0.0131071994578363, -0.273621154418411,
  -1.05187304113107, -0.690792351201063, -0.310145251722981,
  -0.419232391022748, 0.00207848010512483, -0.322282419669117,
  -0.0496906281799162, -0.0568781599424564, -0.136925886672262,
  0.70487089665764, -0.146196572444711, -1.10355818149705,
  -1.08155901610402, 0.465033266645263, 1.30720555196323,
  -0.168866031764653, -0.170478254633812, 0.194726706323857,
  -0.189176878182768, -0.111883222854729, 0.664624202707357,
  0.168244277753026, 0.119010173285873, 0.0169634768614554,
  -0.113346140480676, -0.0855363062971433, -0.0349556652336281,
  -0.0513204237882002, 0.0135891866341755, 0.895107954732681,
  0.638262300191758, 0.228255814448113, -0.438738504450138,
  -0.387010922308603, -0.100716607582027, 0.00465774588774593,
  -0.407785614715242, -0.0322299875750706, 0.372025272091921,
  -0.170250848543308, 0.058225974732947, 1.24809969265263,
  -0.0231762297016824, -0.194781585127138, 0.236236092214142,
  -0.556378351959913, -0.24960624988394, 0.428999562435163,
  0.0562585903465788, 0.274829648174137, -0.618012101754937,
  0.22960006361401, -0.397985448908625, 0.224341785611677,
  0.242383663637778, -0.738284461835436, 0.0638402842234033,
  -0.0427334618456871, 0.0770288148881546, 0.028989568676523,
  -0.0860381741856761, 0.229788952053054, 0.238801611395318,
  -0.0637731635771994, -1.02441487412722, -0.167008035286386,
  1.25088952944505, -0.141641570365527, 0.206644179022605,
  -0.00371192003273734, 0.322995237772875, -0.202671166349023,
  -0.717872729221864, 0.255199470323838, -0.539472111739068,
  -0.845133195889184, 0.139190109215433, -0.472115801503397,
  -0.193504178140171, 0.184608920960382, -0.145297294533941,
  -0.558330522842037, 1.3284791559216, 0.0263512192849006,
  0.542058657756367, 0.98737068944574, -0.0316313947323882,
  0.360044098655504, -0.0307720186991017, -0.169172839697253,
  -0.158326730783156, -0.683299038830812, 0.547849756298512,
  0.376380179147994, 0.304637519724526, -1.06157902829186,
  0.318969504881595, 0.0113741889096466, -0.171589624142154,
  0.315056778565434, -0.0325993044759429, -0.565169847170513,
  0.510017971715141, 0.408224521103148, 0.0334301567058064,
  0.209374528930822, -0.0344607681520465, -0.434613462181884,
  0.204326366835063, 0.155148624612996, -0.496470326069708,
  0.178803604647801, 0.275905242176702, -0.0143458781248039,
  0.471341158710422, -0.212320571402324, -0.116888369935281,
  1.13163177516956, -0.401744304102691, -0.0595470214296693,
  0.0406409352066271, -0.719991103227649, -0.0304720731126693,
  -0.0493063512400351, 0.539573471678809, 0.366666261601722,
  -0.220124571791151, 0.429972199832907, 0.312621762079206,
  -0.314189292894685, -1.08800901959671, -0.227233874404022,
  0.324497788109461, 0.160014567478713, 0.24840560700296,
  0.272529476538695, -0.082230098200535, -0.402308265712138,
  0.337661563734205, 0.408730836010278, -0.0654484535005315,
  -0.117426517689273, 0.18530935544306, -0.233376557077399,
  -0.397782501765106, -0.226245552249892, 0.580562787244865,
  1.71920231803835, 0.951938073820777, -0.414391004974177,
  0.836920883383325, -0.415262896584956, 0.0218739778684719,
  1.0242121167373, -1.6510852884564, 0.933962565404589,
  0.873230228404082, -1.06020907816404, 0.377702457017104,
  0.220410034260708, 0.120408286908575, 0.146897075428373,
  -0.233389884907084, -0.160256717852732, 0.0789140827357768,
  0.714091761279033, -0.276877406737522, 0.0417942177063557,
  0.289353528128453, -0.0369116513785321, 0.0795743085285621,
  -0.0397045887475011, -0.18844801156417, 0.272149009983669,
  -0.242964898517945, 0.262315439887467, 0.415461987316961,
  -0.141675787529418, 0.246076477959494, -0.168297390607416,
  -0.357317842416117, -0.328294705914413, -0.64733143474038,
  -0.116791095930639, 0.23187626816048, -0.800432666695531,
  -0.0497978548951061, -0.279938171796347, 0.323566334573361,
  -0.812036899321848, -0.794780657486609, -0.51072600415361,
  -0.285507030625019, 0.512483504109157, 0.477032000865849,
  -0.0277766042147359, 0.17449949985163, 0.0976211989740954,
  0.112656446984609, 0.370324554896839, -0.134819628665873,
  -0.565188473086988, -0.354743662375693, 0.781688850328131,
  0.253366770075377, -0.133114200318179, 0.0524429620281874,
  -0.276825746829871, -0.858777940164077, -0.138928163854005,
  -0.281450718203631, -1.37102582293886, -0.511834800050632,
  0.182265478633279, -0.222973774668573, 0.101940043009118,
  -0.649590096090393, 0.667883622240404, 0.401384787440746,
  0.618877416099573, -0.580332681086581, -0.0348645263109774,
  0.297871577779791, 0.175708180676272, -0.115751039314497,
  -0.289195286788445, -0.284448484320039, -1.4326832083921,
  -0.588257797722855, -0.212942604170061, 0.62980599004536,
  0.14522515006445, -0.338416718453347, -0.0719811970403851,
  0.230311604809338, -0.378477394006534, -0.423423603613413,
  0.272470632874817, 0.712316594651635, 0.468322329312266,
  -0.0249661560542972, -0.0227570511643196, 0.289907876351478,
  0.0953424836664244, 0.324900280585009, 0.0374881162456714,
  0.35884328168174, -0.289558676974222, 0.0585722620440683,
  0.122745133226602, 0.100057547239726, -0.195936422918073,
  0.0644112825320025, -0.210054692483299, 0.429514093444298,
  0.34714264745814, -0.0146076376056645, -0.295024110183377,
  -0.264405825422883, 0.0834882759341405, 0.0795686400968585,
  0.133141680988093, -0.161036730951586, 0.0800614507437729,
  -0.464545503956033, 0.627782776176712, 0.302988081283066,
  -0.336281904377697, -0.0144582695881471, 0.00164690868470343,
  -0.218920818993404, -0.180723167888098, 1.27039564691362,
  -0.813996211245982, 0.480570879848237, -0.410011308167146,
  -0.30313373651757, -0.184795066950793, 0.198105085029584,
  0.658570995004448, -0.195113942282748, 0.430478366194183,
  -0.84184597744434, 0.128979296104243, 0.230929844730867,
  -0.188634557492053, 0.0162861317211379, 0.105941730179998,
  0.00810969663589278, 0.0187010780024251, -0.0239216567274075,
  -0.651793367502972, 0.340607924981084, -0.0633647365934914,
  0.103603976616134, -0.101096720445605, -0.293800702707223,
  -1.59143699627703, -0.463444852485517, -0.275008499951014,
  0.188681058053373, 1.11125201548625, -1.88549552691266,
  0.283228344628538, 0.0413860510875813, 0.191360524365733,
  0.249846437557075, -0.080432718523442, 0.268009999565841,
  -0.0999142532201033, 0.763687223796392, -0.234595556763957,
  0.0901411612013329, -0.496173647677684, -0.0343980993580323,
  -0.83805639541887, -0.400331870298174, 0.339301949254142,
  0.229554992342924, -0.930892952503313, -0.76665634209746,
  0.278870597129073, -0.0294573877845954, 0.189431208745321,
  0.250231995256229, -0.343428338572952, -2.28037640757929,
  0.370491074092436, 0.0794657822320328, 0.175025315286084,
  -0.161879143037084, -0.00629986204280725, 0.130257953093848,
  -0.467363428485739, 0.760108541753219, 0.285504769509169,
  -0.298182014173816, 0.246900048493994, 0.188282937302818,
  0.145783456876764, -0.0481619329646669, 0.0161143057491261,
  -0.0504584986534748, 0.078444229283757, -0.746994115096354,
  -0.204382710719975, 0.337528011555356, -0.610720150813078,
  0.0301342943379586, -0.202696759766628, 0.117823054361133,
  1.20957783517611, 0.849099735380018, -0.629099618611954,
  0.821250314455495, -0.667408480848148, -0.138026370130076,
  -0.512568564668704, 0.147862942142894, -0.108572217244128,
  -0.543212868370717, 0.101701612782243, -0.478417053226069,
  -0.475898756861702, 0.10969171337381, -0.246952459095516,
  -0.0824910004864428, -0.125722065055674, -0.1647079562162,
  -0.517499490991674, -0.152344005492798, 0.0652597460594407,
  -0.686864677156272, -0.260234218515415, -0.559053239954506,
  -0.213430987568739, -0.450126390856665, 0.0795656535691979,
  0.242161039548692, -0.508837686956215, 0.113298739585723,
  -0.135490377467353, -0.41659766428283, -0.085529170249319,
  0.0486867183941303, 0.0840984126555795, 0.351967033340869,
  0.618344531450669, 0.153660857494661, 0.304118212638999,
  -0.0475165203732438, 0.306577779964178, 0.307712184066683,
  -0.138349560463867, -0.435451908513439, -0.142590479748829,
  -0.157180703848283, 4.01988605308068e-05, -0.309263074994985,
  0.836009120539432, 0.922138474233192, -0.140827135533428,
  -0.00961580154267039, 0.366281301142221, -0.103495810850569,
  -0.563747850355421, 0.493846801385625, -0.678254878911888,
  -0.715576888312091, -0.150631855330234, 0.00446219250860145,
  -0.0712419306041977, -0.0491533178322363, -0.181481388592094,
  -0.117463153272034, -0.25577441872639, -0.0235361429370499,
  0.504836308027494, 0.391817275697362, -0.181597773496231,
  0.166774123576601, -0.156849405722187, -0.508300300769258,
  0.21467435310833, -0.0917601588536223, -0.142507377190615,
  -0.181516595932459, -0.211063158584257, -0.665207659916138,
  0.222179306332853, -0.104242918966565, 0.277512747917031,
  1.95848642932234, -0.517139904520447, 0.527619341023627,
  -0.691299273429573, 0.230294207366673, 0.201453674495634,
  0.0568611314587897, 0.200818099462503, -0.0454357798796376,
  0.652090660170742, 0.15211809080501, 0.626706155622609,
  0.351351877402252, -0.185005266041323, 0.256550968075215,
  0.423740900285307, -0.0741867887093387, 0.0667073963384699,
  0.380116621149999, -0.0598780727782894, -0.185606253964907,
  0.604256225950872, -0.0407169364656139, -0.649252809377556,
  -0.106287479307992, 0.125106387766443, 0.294443216599934,
  1.04857923489436, -1.41002656614875, 0.530763844551404,
  -0.421613599293166, -0.777079400828128, 0.766877623491602,
  -0.0891793761376393, -0.161907714785229, 0.350797688389172,
  -1.08228145431118, -0.320494516880555, 0.996793581949202,
  0.845266746473958, -0.132889778475034, 1.13065920611296,
  0.0999297323594728, 0.0214089018000361, 0.178797351594005,
  0.449289218188335, -0.246966730431642, 0.220635369788342,
  -0.463279110702699, 0.62711435097338, 0.2864023130374,
  0.35989592080089, 0.243143796024439, 0.262883417144296,
  0.0934262620781316, 0.241083490451358, -0.0554265517486415,
  0.136793651816458, 0.041837299148189, -0.658663769605551,
  0.133372486605705, -0.0977655979346535, -0.0854273469645034,
  0.188114701328114, -0.259721459341595, -0.00217030081237521,
  -0.284894035221984, -0.745275717595078, -0.145715776656184,
  -0.16406478908652, -0.0958820731979478, 0.0378509734650617,
  1.29411973502747, -1.03143477338246, 0.195653934576503,
  -1.04708552883484, -0.289622889612558, 0.0320639514709839,
  0.257108049634739, -0.139624405670285, 0.0276098065322393,
  0.189683802317638, 0.259431768997604, 0.888230541482439,
  0.484814334214337, -0.132820956342153, 0.154706625800596,
  0.233818757390063, 0.239075852783807, -0.0588586690286524,
  0.875446573442691, -0.281046849196777, 0.0175399220246246,
  -0.347612329187386, -0.270009838318105, -0.410151800921706,
  -0.0574413060344248, -0.0117053838059625, 0.0623585253843607,
  0.118691129463468, -0.103637029574337, 0.52574488208345,
  -0.0927957533638577, -0.633150107911917, -0.637547437480783,
  -0.0915282011169298, -0.531098945349423, 0.168947988282132,
  -0.946733685448669, 0.320258976255044, -0.400856146027943,
  0.130841231889968, -0.668787213667241, 0.574795428366866,
  -0.346603135546072, -0.268642492632926, 0.29658033687634,
  -0.435915397303957, -0.368850360402146, -0.675781383473421,
  -0.587046677590869, -0.621677442754282, -1.78004053394199,
  0.0890305662772982, 0.0360416192426774, 0.203738110286824,
  -0.196170997554309, 0.425374979393467, 0.110994327760366,
  -0.0503619018245659, -0.265620418842201, 0.0390500727458771,
  -0.412805976017877, -0.133094356179665, -0.120581240567986,
  0.227705525402635, 0.983386007654127, -0.661088541676972,
  0.516375150849937, -1.12967229923081, 0.12219025130904,
  0.00831289234436075, 0.365502339522865, 0.0230628448190919,
  -0.0598082042673235, 0.193984911992983, -0.124668583637525,
  0.0332518780693564, -0.167841700651835, 0.0625105856107012,
  -0.38553933332714, 0.0106587144551577, 0.047690365347055,
  -0.453893971862764, 0.240073438421142, 0.0657280319231405,
  -0.211563614900879, -0.0171567354373214, -0.239717827117181,
  0.0237414238036049, -0.325290572829616, 0.186200329411783,
  0.144683522976166, -0.28553653513078, -0.152913775979381,
  0.29386075444972, -0.6790014706374, 0.0501027692214804,
  0.0568309242169052, 0.0423299027384605, 0.185273227636787,
  0.0379245485103113, 0.30041483303796, -0.486701458554463,
  0.349451701895569, 0.354628741849918, -1.15233829265583,
  0.129236325085095, 0.336136928043264, -0.0563151703717112,
  0.191687723769609, 0.278552162992804, -0.0493500564444272,
  0.197964379172471, 0.283666477247737, -0.0810233613067516,
  0.0817181369790156, 0.140618362666475, 0.05441568061406,
  0.475465003684118, 0.123837218934749, 0.442841634452316,
  0.395455474654944, -0.685858420271735, 0.181398766409053,
  -0.293846413412191, 0.18534077729579, -0.0596831308389717,
  -0.163357158275428, -0.339591380474217, -0.477329672753629,
  -0.28409682211495, -0.114918980498397, -0.310798846897346,
  0.0907670027629759, 0.0356492067603759, 0.345149148575281,
  0.501809399127437, 0.525488216667568, 0.0277930138709548,
  -0.949349889172347, -0.551102258583743, 0.638462434304533,
  -0.144386784349405, 0.0478107548779532, -0.0487028738190789,
  -0.269288705567351, -0.437710286912995, -0.491761368484878,
  -0.29240002471729, 0.248182395355864, 0.101006870593198,
  0.198477421100009, -0.216294228086155, 0.0143832302903482,
  -0.40346790792497, -0.339117819701558, 0.0804123901991985,
  0.115108418662002, 0.38876464774225, 0.368626574073217,
  0.279243664062168, 0.190843275077013, -0.322082102468966,
  0.557546499967885, 0.110715337846471, -1.00979877753078,
  0.705773152344735, 0.540825102258059, 0.0881323704986467,
  0.128533713896126, 0.301951388921951, 0.169142466955922,
  0.697849048213329, -0.268618058077957, 0.378666097934881,
  -0.651732636887346, 0.738667452113674, -0.508329588606488,
  0.340367374053484, 0.200271899919297, -0.0823367313910278,
  -0.401444374592157, 0.161564443454381, 0.327458051990912,
  0.936964184286183, -0.237621889986319, 0.0895158818485099,
  0.132766420039099, -0.0515261755197276, 0.31285279656253,
  0.175605332878886, -0.438192561257727, 0.226092498095669,
  -0.348238692061781, 0.767242383530324, 0.620219883704266,
  0.247142066005552, 0.163014665021789, 0.131462540620302,
  0.159110595811905, 0.135819092633785, -0.0756124700588107,
  0.32673762567934, 0.0825993811862784, 0.777870717464528,
  -0.370887962283647, -0.236065631722922, -0.194928901195106,
  1.72201261082371, 0.00947019751309562, -0.347563906265374,
  0.0680470695146651, 0.0191757552007686, -0.328380189008071,
  -0.261083845747734, 0.00845243205905241, 0.0353631320009814,
  0.14717378847342, -0.238514871637136, 0.319011181413703,
  1.10909208618213, -0.703758559570137, -0.0435145036207595,
  -0.211116327982721, 0.156706023517194, -0.300268107871057,
  -0.564905090454177, -0.116633207169653, -0.543121751303117,
  -0.818585843513278, 0.397329377222964, -0.612681354839417,
  0.017812014521462, -0.0346184780640765, 0.0082174513226979,
  0.295132484413035, -0.40054152659519, 0.156146143225882,
  -1.68040080802289, 0.987415280990581, -0.418842654824823,
  -0.259717621181266, 0.0809608981281909, 0.344762987850959,
  -0.942474018067098, 0.0409431546460739, 0.745447294999559,
  -1.58579273475185, -0.583708847455147, 0.985394066839514,
  0.258912744782248, -0.0989703255550896, 0.209238500696728,
  -0.169222335822336, -0.223235175887048, 1.22812608530356,
  -0.664198644496171, -0.275675183775019, -1.02215101435919,
  0.185762874645491, 0.0652106663358479, 0.0436960141514642,
  -0.696081342236382, 0.657961172425268, -0.0590068609040234,
  -0.0939905420828469, 0.31812283742504, -0.00172050579394634,
  0.307578765053199, 0.0393493342342992, -0.115406662234474,
  -0.552274110002296, -0.188043520379149, 0.253504478773653,
  0.195303606996157, -0.0537472371423025, -0.107140319990729,
  0.169919714542381, -0.109611840179161, 0.0887740670949165,
  -1.39380644568458, 0.439293663997803, 0.569826564500841,
  0.0679688409715019, -0.415300781999993, 0.0686627818020778,
  -0.1340128587755, -0.0395410374789246, -0.180649866177488,
  -0.221273473979366, -0.0229636451244886, 0.126033300083321,
  -0.30044731198421, -0.11001408341098, -0.0624326275566202,
  0.26093022532863, 0.078869768673072, 0.336467551260967,
  -0.0599838707061267, -0.180180665987926, 0.250153134087915,
  0.0735399395498073, 0.310289317100224, 0.393163714507256,
  -0.156976655726957, -0.0711648288938424, -0.0420898121846291,
  0.0646759519492794, -0.403884973948937, -0.252927438649135,
  -0.0198460931691664, 0.93407474261077, -1.0146879998174,
  -0.302093100912614, -0.216251105633622, -0.365334857423843,
  0.00617436872720658, 0.101710359985308, -0.379160419403031,
  -0.163077791858468, 0.280337283007175, -0.7316568264805,
  0.074026112603745, 0.0521762064321673, 0.0677921747870854,
  0.195985418347824, 0.454965194163611, -0.63666195851072,
  -0.340904333112812, -0.106509061623518, -0.228974827758092,
  0.208318305028826, -0.0954737777826645, -0.101821649348041,
  0.72213680559536, -0.652888506805695, -0.496595236601579,
  -0.819797263581684, -0.474972358932433, -0.0773596158621223,
  -0.264789892696036, 0.0982238158642301, -0.0553096793781458,
  -0.970756089795628, 0.736262900162179, 0.414700666444753,
  -0.108327307827803, -0.531962957345558, 0.551192113463096,
  0.107455954322177, -0.248505402973182, 0.109072086448979,
  0.0499050856641217, -0.0303399093956365, 0.138319222632443,
  0.145885604452862, -0.142125582601298, -0.530514309139391,
  -0.0945166923053331, 0.123476410409976, -0.0202849622168449,
  0.777425868844023, -0.362166845725995, -0.0821498620814418,
  -0.0172452234195961, -0.101267242302291, -0.621618788386041,
  -0.349078641471288, 0.0371389066153071, -0.0509212484113332,
  -0.046642942925161, 0.0232792104936146, -0.185425453179379,
  -0.579245746494036, 0.221395917651016, -0.306744688019485,
  0.0228372512409546, 0.150474110206565, -0.0872799565929347,
  -0.432862775620978, 0.460398055457465, -0.859189622815782,
  0.514309668104127, 0.490855239119491, -0.403010505563415,
  0.240118921881786, -0.00448643990711727, -0.0504151638385455,
  0.281335505835128, -0.00860877678607565, -0.298789810817065,
  -0.0549422134813082, 0.0769193804293865, 0.788718919581685,
  0.20328157442979, -0.191474176578087, -0.276315684153054,
  0.0296520144821887, 0.0411089970630018, -0.45640095238978,
  0.581470003221321, -1.37853348955001, -0.243790002170671,
  -0.279839952773492, 0.135613828087698, 0.098821390273122,
  0.0344843414613523, 0.838561744570938, -1.32972433707187,
  -0.311994025263638, 0.185439646389022, -0.389210295661502,
  -0.185378947456333, 0.0157481144910984, -0.181889475684966,
  0.263237923432507, 0.938534688522058, -0.00070514064902974,
  0.123204625329948, -0.544477712367507, -0.915939319813511,
  0.0108670087997897, -0.0368885971081732, 0.085985071194387,
  -0.781377462193309, 0.439740304286901, 0.416378023704159,
  -0.502650269173444, 0.0195424603686539, -0.0482047870010406,
  -0.139662251428426, -0.124749604975685, 0.0673463176479086,
  -0.623938011653272, -0.226502947474014, -0.62786848657822,
  0.194965642122123, -0.0259657843699103, 0.658136219357821,
  0.0690468130880041, 0.255558863934666, -0.0648812341812541,
  0.624177357141865, -0.376752317340908, -1.31358817720342,
  0.997124512205083, -0.647661570997363, -2.26771004469419,
  0.213866567799588, -0.137151134491985, 0.0865716637776342,
  0.226362356588395, -0.0745121271893711, 0.355263959065708,
  -0.0823298528022676, 0.178833856011984, -0.00808103195037309,
  -0.128061577316108, -0.229885903143378, -0.127781093161712,
  1.3929926658262, -0.0138218123321028, 0.0728226296854477,
  -0.245838399565546, -0.747800972034726, -0.0622479327356794,
  -0.0172058042914862, -0.317349064808566, 0.489658728098709,
  0.822467091239325, -0.659286573854312, 0.427350138521227,
  -0.787362915041189, -0.847164943360718, -0.516795242509964,
  -0.217564801228537, 0.261110146803019, 0.312296902447923,
  0.00551448220685394, -0.809473938529123, -0.0491653078619229,
  0.613198753081455, 0.688025350016965, 0.144225408320007,
  0.285572425957743, -0.0546930869526837, -0.175174286767347,
  0.136894785960099, -0.0243986479049556, -0.0938291074625051,
  0.660637654290532, -0.602954203305991, -0.19060863455661,
  -0.122539317075516, 0.214920901270634, 0.0930336264772913,
  -0.557191370078697, 0.395212355454429, -0.405528650927638,
  0.558275522193443, -0.0761327436071205, 0.844236718385388,
  0.194088955861884, -0.344911306890728, -0.00875017672116731,
  -0.70949379420079, 0.2090482617413, 0.627020575126682,
  -0.790608682948047, 0.345268837489244, 0.433948797538139,
  -0.00957267412519621, 0.152937472283227, -0.061325402188655,
  -0.384019611909548, -0.902251947135081, 0.0698297072558913,
  -0.115270435049804, -0.118259289205182, -0.0693916868299316,
  -0.0109594319092138, 0.137441682192498, 0.024596062553228,
  -0.553020791884355, 0.109995111836306, 0.977719537923639,
  0.2879431945844, 0.963411825364038, -0.729615507743608,
  0.126136655132764, 0.0305995445940964, 0.275358968390769,
  0.692293419641944, 0.515669215108189, 1.36248983132166,
  -0.417797631399914, -0.691884167968524, 0.522266938696197,
  -0.122064073534882, -0.092710775220929, 0.0153263778092249,
  -0.165838534465129, 0.552396026451409, 0.51900382421535,
  -0.116523827218553, -0.81638694741579, -0.443921315818883,
  0.148710986911163, 0.234569127779272, 0.0114905686251366,
  -0.647217967298751, 0.154853724576744, -0.402373785328487,
  -0.28173067059651, -0.0284687101121178, 0.495909830160418,
  -0.0863765203844272, -0.370827074770164, 0.0483744356128617,
  -0.511906546868728, -0.470461418895467, -0.26722680451515,
  0.421536250482521, -0.198460180288292, -0.383206396369653,
  -0.168418054314325, 0.519394829939512, -0.115973783977875,
  -0.858958176640289, 0.317911281629958, -0.39538489678438,
  0.419807402924064, 0.394361534964315, -1.09879256473913,
  0.0463882574181143, 0.374647729010818, -0.189721671805189,
  0.386634276224803, 0.639351921098192, -0.742676494832333,
  4.13342347882761e-05, -0.326335079387692, -0.296578136205124,
  0.338663832619327, -0.00865026456991334, -0.29503107518241,
  -0.20269019438336, 0.0654257941652907, -1.48757724898888,
  0.17087473210553, 0.004229959746886, -0.0488069130822608,
  0.118819546751396, -0.133751360300859, -0.0422437408844381,
  -0.203406317022861, -0.28851203206465, 0.629455097769555,
  0.380668423949243, 0.467865324275709, -0.187518462469486,
  -0.0146619164769233, -0.174346753159202, -0.338156261808763,
  -0.3597696298507, 0.356401560828453, 0.830377714324505,
  0.0548832918348875, -0.471112926373869, -0.307569291705614,
  -0.0283117136852537, -0.0777481171232466, 0.190982033160154,
  0.600489704835588, -0.24535368648667, 0.297880690782688,
  -0.645842102926612, 0.491078762114439, 0.0363426773627661,
  -0.0310044103593233, 0.1888107795885, -0.283351067311006,
  -1.64517539101399, 0.713352149453152, -0.270588620131716,
  0.351861491194999, -0.302748478625049, 0.324987735004108,
  0.289239219406916, 0.00962225204675738, 0.253307630945086,
  -1.03453893021987, 0.0682504850354597, 0.502085917305878,
  0.372708354335114, -0.0139743235386671, 0.524978983789687,
  -0.162612177866715, 0.247589559143759, 0.0274339508490366,
  -0.0130371299065236, 0.228213877542561, 0.495229106030191,
  0.269421045996153, 0.277776090332224, 0.566183573979302,
  -0.0555194385855366, 0.00115428067923005, -0.34182950533502,
  -0.25144932895663, 0.130375730093625, -0.170138949149915,
  -0.214883312301113, -0.347894750169904, -0.78073759016473,
  -0.053475363420489, -0.233892548063756, 0.235995802221291,
  0.120224741144865, 0.590181481541618, 1.20820053202953,
  -0.0255235070897534, 0.288649158301749, 0.87438895494921,
  -0.0815036580797776, 0.199353831147257, 0.0581278037938487,
  -0.116810287708343, -0.30964988633057, 0.423992997518599,
  -0.2338811502123, 0.804353377388209, 0.375466042767789,
  -0.0420917498048826, -0.147583991209068, 0.332046847650128,
  -1.44640931907899, 1.37149074696574, 0.60680893571311,
  0.474702200843643, -0.787313672350555, -0.18206592306842,
  0.156843464978844, -0.0928150591605268, -0.15098408905723,
  0.116695990410461, -0.75297073244972, -1.80110730861946,
  1.24909651391949, -0.0827025135298681, 0.134437396554048,
  0.289844767365687, -0.112007022418903, 0.0196901918914781,
  0.0103604028332825, 0.0709398185042936, -0.0531379348096264,
  0.849075607503787, -0.836468998578208, 0.256302733443072,
  0.177337316285967, 0.247834658920927, 0.149388015251655,
  -0.0376220947800356, -0.229783100792678, -1.45858201920388,
  0.720651895947477, -0.201627766477682, 0.074859736756434,
  0.0929251166754792, -0.232788182288144, -0.359334603736239,
  0.226081085794195, 0.988805191370781, 0.22921093672956,
  -0.683048585887352, -0.349958438704557, -0.859886468330819,
  0.283642184837268, 0.325265525217744, -0.175292779384396,
  -1.06650928764236, -0.0488533344370842, -1.2237942340614,
  0.493136827934238, -0.0116613193675068, 0.883546776412794,
  0.0218878964214764, -0.196533877244895, 0.341047216599913,
  0.963637420051237, -0.568670211641046, -0.616752617468845,
  -0.22998169874762, -0.00282970701808322, 0.586610619490287,
  0.330489586948142, 0.21449788224097, -0.108246936892692,
  0.0851040917896065, 0.193616957818985, 0.378371131659755,
  -0.254690259931135, -0.135139578946369, -0.574266752257138,
  -0.159351039930394, 0.20677123512792, 0.00800400457562319,
  -0.218760404883293, 0.250339511401248, -0.472231217893496,
  -0.0821757687373654, 0.111963389321754, 0.0713664520724097,
  -0.0232743145168702, 0.213485117671828, -0.232006972098378,
  0.00473088768624929, 0.240738148122606, -0.113713113002847,
  -0.147232167253857, -0.0485904655112181, -0.88183667627805,
  -0.187065498650166, 0.214409517047549, -0.108585963067293,
  1.01432690438985, -0.000303315356698167, 0.250595659322862,
  0.564011393710354, -0.243840974917496, -0.50620466338044,
  0.181973939938499, -0.0313137844699003, -0.40118089241181,
  -0.246959919390946, -0.0709441375305839, -0.803333681041228,
  -0.0726034543457055, -0.471254080942975, -0.220801182738676,
  -0.03506528890436, 0.32076924895169, -0.0438299535649884,
  -0.739771030725519, -0.14788656099402, -0.667449281597168,
  0.484976545061237, 0.0636126606785121, 0.124794815664252,
  0.217700409998173, -0.322703229143718, -0.167999046925187,
  0.21653691984845, -0.360141530299983, -0.123717112123872,
  0.0856101167415886, 0.236195720580547, 0.169102275394217,
  0.0630909646763585, -0.181673450287553, 0.19354038674415,
  0.452686259850985, 0.0223398677567956, -0.129371697969697,
  -1.16866636720383, 0.417897457456154, 0.734605568960296,
  0.0590496712779499, 0.0215479197616641, -0.218472612734029,
  0.350304686157352, 0.0489222310939746, -0.865244880178951,
  1.45761898559072, -0.63329654000341, 0.207345189258054,
  -0.0516509829964578, 0.0304421329221757, 0.0100862871030431,
  -0.328643856269061, -0.612328765394685, -1.41014910319772,
  -0.244375674296118, 0.536566500788029, -0.804566145490398,
  0.124814782753675, -0.173871110468016, -0.36664893667458,
  0.281903448674142, 0.0564529515451286, 0.825008812180433,
  -0.118495335225794, -0.777364074035202, 0.413834099669893,
  -0.0727651524836561, -0.388824276770612, -0.267658608945131,
  0.0602658313188705, -0.0739902789353298, -0.206765348994904,
  0.181797273544619, -0.621315135884717, -0.299900537109158,
  0.0924855323303687, 0.298785264863642, 0.0640128081934286,
  -0.00282319565256329, 0.55716838255747, -0.188970074395083,
  0.110313320398009, 0.0735054274874937, 0.274282407354477,
  -0.175965443383218, 0.218194642792508, -0.000563044109719954,
  0.0831140667743245, 1.28621728342335, 0.685418727041812,
  -0.948735628739112, -0.14436544873674, -0.677522211683737,
  0.487374337619383, -0.22242365483448, 0.0371339889999224,
  0.607551737975646, -0.0738685947711644, -0.0677397737258717,
  0.623044679842183, -0.0660868993867115, -0.191382492387963,
  -0.100995215231051, 0.14790018752512, 0.0291269246664473,
  0.332899596508221, -0.0673387902687161, 0.589506082414742,
  0.32108022085013, -0.348628279516004, 0.642544949061282,
  0.204488887786842, -0.0108483664528518, 0.332155050703468,
  0.0120742540278173, -1.3603020763889, 1.81032730693711,
  0.0119005218754614, -0.919285496428318, 1.48495336441012,
  0.0353284338520237, -0.149226847651338, -0.315233532348949,
  1.02135554704015, 0.339915308681229, -1.02134621596716,
  -0.438028744425051, -0.101993763235886, -0.587722876342148,
  -0.171504892748695, -0.0118663982456807, 0.299897127709396,
  -1.08679582371284, 0.451099940584943, -0.467793363359806,
  -0.661084371229145, -0.646159284510926, 0.472118406375993,
  0.234308196158552, 0.252022077704367, -0.150060490114457,
  -0.373330176297622, 0.724776669303702, -0.856597655022632,
  0.187336678932535, 0.211114418994769, -0.273436542945818,
  -0.242663558363736, 0.225193460723068, -0.0942705230078985,
  -0.0325326529522282, -0.582941914815521, 0.382779387622727,
  0.275857076295717, 0.391779935174511, -1.28959362740954,
  0.0234900013744077, 0.281547638397373, 0.0428759720107508,
  -0.36873973362301, -1.04007294534848, 0.224350776097276,
  -0.395346946571072, -1.64146252289358, -0.000728370511095287,
  -0.0528517709808298, -0.149042527137762, -0.229979586156217,
  -0.187013758728473, 0.254472519461497, 0.701061311211169,
  -0.580095561853736, -0.608956791342806, 0.109256939365418,
  0.161063359971421, -0.126056563417316, -0.127028977822747,
  0.0309295804326417, 0.466962436044629, -0.00509902293097431,
  -0.0144001999530693, -0.891424874570547, 0.0453201092448083,
  0.160107289154327, -0.00656365711484253, 0.0757258112847941,
  0.366295391088042, 0.718132292883207, -0.35276581230663,
  -0.756562126884579, -0.886775466919, 0.39444677773146,
  -0.0681569520874959, -0.115725370542541, -0.11064843401706,
  0.714016793784153, -1.21295400552144, 0.136068349568972,
  -0.532766241660877, -0.686893841236032, -0.00563356507866633,
  0.195528470117995, -0.268883976216776, 0.04283968786927,
  -1.03953380284929, 0.108877317682786, 0.553392662976291,
  0.888143830703823, 0.849813244769084, 0.268314582112027,
  -0.0377072794061449, -0.049552037273404, 0.0468431709865009,
  1.40973325355937, -0.0646770949125015, 0.863288954515979,
  0.77487147181165, -0.341230411832046, 0.0516023353675032,
  0.147082077897471, -0.351943557723487, -0.0771874746747209,
  0.143275340690474, -0.314624723956782, 0.0174450869705152,
  0.467513481899318, -0.646702131858923, -0.285270922288497,
  -0.179543510741771, 0.0858664473339743, -0.447741691040381,
  -0.29358268840547, 0.0283341661008289, -0.419173906558653,
  -0.154315285016607, 0.249615282429677, -0.416723568617703,
  -0.142945959783797, 0.0440690695265452, 0.0893239667587201,
  -0.112570979014603, 0.357824830609688, 0.371829689760982,
  0.389944985271175, -0.23931361973022, 0.100038973276065,
  -0.106074690849474, -0.326457307289432, -0.112387725689739,
  0.492176219622584, -0.378463387480207, 0.352473319410793,
  0.231584432860482, -0.275915293409337, -1.00029541541031,
  -0.156664317284257, 0.0967056529489213, -0.164028031245945,
  1.11176772493685, 0.500474609204391, 0.0490269618905728,
  0.744493772261988, -0.866383666069416, -0.576440591024884,
  -0.0371576507132238, 0.123086354443483, -0.159366253522306,
  -0.170852160314503, -0.547668511879002, -0.0736187043377147,
  0.204819395671962, -0.300410969600196, 0.36019380696446,
  -0.0211896304622535, 0.410069668019505, -0.169479745975584,
  0.293414914858135, -1.16101087215201, 0.0480994235404731,
  0.156779253539235, -0.479958170930831, -0.0427530662549751,
  -0.0175494452784145, 0.123607084297787, 0.147273326087932,
  0.709505053751468, -1.05108843750475, 1.40826650903127,
  0.64288493118134, -1.00666081122908, 1.29955929572032,
  -0.0806677416788809, 0.13233330115143, -0.00686706597990262,
  -0.406933117456058, 0.202464641983354, 0.373528725720593,
  0.144081208228742, 0.039286127837329, 1.13595937514716,
  -0.258221881722504, 0.27775136982805, -0.240934301444888,
  -0.428429984632277, -0.89567118899695, -0.873063017051456,
  0.721861258392499, -0.037431713222883, 0.220607855709633,
  -0.143605973719434, -0.288070459800507, 0.344905456065778,
  -1.73195998850439, 0.480039901585336, -0.181991296544453,
  -1.07257250334165, 0.965296449629971, -0.022691778063617,
  0.00156901228188503, 0.160835699310354, 0.133340979613421,
  0.446280512808721, -0.141027353702054, -1.11420335944111,
  -0.496643716164842, -1.07727591361375, 0.194860531971344,
  0.141361514152254, -0.087777352073299, -0.0353328504258796,
  -0.260997085426142, 0.656144767209204, 0.906308123166132,
  -0.0521789402846826, 0.164407672673971, 0.0548651736863894,
  0.00523972737299356, -0.228894076078977, 0.259591281314655,
  -0.159578181556275, 0.750372961595211, 0.606722401649977,
  0.41945339640432, 0.523687855604783, 0.201327017812372,
  -0.0220672727451084, -0.0639132118280522, -0.0274584562601919,
  0.139081269697606, 1.15133467935976, -0.40621169039793,
  -0.240723343958671, -0.0145550221693133, -0.438789721616196,
  0.28793337484176, 0.0740038493568701, -0.123840377369809,
  1.06632718800203, 0.859184388596857, 0.490203580376076,
  0.259511188175147, -0.0808602365901273, -0.533244933291745,
  -0.116440780378283, -0.162489042073293, -0.233012727406893,
  -0.238961968536958, -0.512096334281456, -0.271452730121786,
  0.0913580295629367, 0.112277070424457, 0.0831573603841146,
  -0.0223089847485181, -0.228180789967761, -0.131514094474195,
  -0.17927139363527, -0.4374499823399, -0.041443751082297,
  -0.030242357119724, -0.244766148103739, -0.376207089112575,
  -0.193941373453969, 0.0324751182624099, -0.023304101676328,
  -0.385402528587496, -0.0103519547679927, -0.14685624908262,
  -0.635388308350478, 0.672100218961425, -0.342400814986391,
  0.050440163873245, 0.192467902675981, -0.092302907633049,
  0.44213449066052, 0.168832029895036, 1.26189046415781,
  0.19712348051113, 0.248733835854212, 0.351698763321747,
  -0.174308796419731, -0.265727802326906, -0.0785372380034379,
  0.647163132196055, -0.449660472678024, -0.402855996190227,
  -0.0855667984414046, -0.218053256298806, 0.603833510011974,
  -0.13400122213461, -0.298194525725066, 0.31454312711129,
  -0.154940179114024, -0.368487510425697, 0.518350892771269,
  -0.0148339656489101, -0.275966903790457, -0.646693764238694,
  -0.256380385422055, 0.200879139068997, -0.181139243601398,
  -0.282415365503979, -0.140866388015515, -1.24277023164821,
  0.160854883377688, -0.224761094639927, -0.351518968648754,
  -0.0560818186156502, -0.388457431749004, 0.0878261997465043,
  0.212295569846063, 0.602987412194803, -0.304259203253538,
  -0.107665959440847, -0.634093525694954, 0.791521517157084,
  -0.250404649481538, 0.0116354777937633, 0.190668172318788,
  1.58210436669047, 0.00738285582135487, -0.155940229161017,
  -0.351996667972628, 0.0105688924761388, 0.219880982158371,
  0.170262380976352, -0.17721444817897, 0.0721379754389649,
  0.558510815761977, -0.792463482014919, -0.38064738704659,
  -0.530614063715679, -0.6600975631075, 0.474131699471196,
  -0.182256379663732, -0.150276481226576, -0.0984784831818344,
  -1.32951266285728, -0.226205943780987, -0.246167789707727,
  0.0419487005466511, -0.609226492137771, 0.288868748562844,
  0.0726158804053857, 0.0817468379675201, -0.110024249814498,
  -0.364727096094947, 0.115103440538111, 0.198555592099023,
  0.486924255246827, 0.429489507539297, 0.227977083465821,
  0.182799347592705, 0.120512332917831, -0.170368804615139,
  1.10754322879031, -1.36068232228328, -0.425013625710354,
  0.0894152674589775, 0.538739005121867, 1.40637711940291,
  -0.041276144853925, 0.0209047094643854, -0.0507062023539657,
  0.352698243954153, -1.63461401807914, -0.0664447196464586,
  0.55921331800135, -0.507841881219836, -0.43014902244632,
  -0.0639271186129423, -0.142492476399077, 0.174889629356778,
  -0.271034455517925, -0.225599322397568, 0.514232037593053,
  0.0456245003146636, -0.449947067524133, 0.042833533339493,
  -0.23851649635159, 0.0904148889870491, 0.0249866607039498,
  0.498891025771626, 0.105107978399391, -1.20316915750997,
  -0.0706210612546641, 0.403917347300564, -0.71525526640608,
  0.0582469162278689, -0.0502112995935567, -0.162385543408428,
  0.51135629564276, 0.342613409689122, 1.89855626936106,
  0.336933748983724, -0.354773849269803, 0.189690749172213,
  0.253015039548677, -0.21347203632479, 0.311685345056292,
  0.243051602263234, 0.0116243392544532, 0.268699787883585,
  -0.110599547906376, 0.61200566439002, -0.199813616397473,
  0.216511644442053, -0.245288626546574, 0.350430696122302,
  0.481988180852517, -2.42785383040832, 1.33413782069176,
  0.617705197595945, 0.981392900333544, 0.189663941226393,
  -0.171605543102071, -0.0965880380294174, -0.0330518044636983,
  -0.407947297942824, 0.17396502174601, -0.186333604322128,
  0.512992508393903, -0.279078897473341, -0.139438696370477,
  -0.219624154098371, 0.0756243323356577, 0.0632476007365198,
  -0.417063390401648, 0.0749436280278535, 0.123814719285347,
  0.361411743458419, -0.294355855946857, -0.120690988468023,
  -0.180818215126577, 0.120297689347579, 0.0497866631637219,
  -0.24733714651373, 0.362409087153, -0.094735414701176,
  0.0664538646536523, 0.424699677162205, 0.196557035423255,
  0.0687719754591545, -0.0352882389067727, -0.171803127248763,
  0.364834171866004, -0.294354197011764, -0.277221205387301,
  -0.259007675443348, -0.0160794820762202, -0.136573158167838,
  -0.32639981112235, 0.0632815084040787, -0.0837348195881625,
  -0.390266694786663, -0.00599161843151497, -0.154612167217768,
  0.168327398385834, -0.29253059969585, -0.33737008763006,
  0.127483520630247, 0.289102945609705, -0.403951829934189,
  -0.182921939537308, 0.174879116675529, 1.34361881522703,
  -0.0324443808457457, 0.522666235202016, 0.570972321956303,
  0.109616521703934, -0.212912913564087, -0.13760244577014,
  -0.192110250041793, -1.49820212016527, -1.46838445498668,
  -0.194470308448765, 0.135422481934349, -0.276200933001167,
  0.0302356421976484, -0.138973691311048, -0.0705672931561217,
  -0.719282227573907, -0.167360802515758, 0.456519967863114,
  -0.629437185553094, -0.185492546153886, -0.0922205876896344,
  -0.20273238876669, -0.384883605382853, -0.416766901409818,
  -0.0891065378449645, -0.387456661163169, -0.265124298066722,
  -0.316150159256214, -0.542793672062361, -0.575948256015381,
  -0.193282690221598, -0.0521323941455893, 0.289490706937746,
  -0.37215408607611, -0.676381959926544, 0.0317440697374541,
  -0.542844410474067, 0.636992305818783, 0.303089423599749,
  0.171746602885388, 0.167415811392757, 0.359775517230303,
  0.630117335926097, 0.0425669023633071, 0.319666824839443,
  0.157653998391078, -0.555883569948587, -0.00217134424968005,
  0.133037412946064, 0.381458069076279, 0.263467062765529,
  0.192396973579636, 0.543539485781343, 0.90976473444033,
  0.0896918432262688, 0.211130937807616, -0.724081675587566,
  0.115613032824522, -0.0262801731124844, 0.106947970010922,
  -0.796898018644467, 0.296127223460506, 0.314424277207787,
  0.243987989112659, 0.550265326211466, -0.785905684607331,
  0.0441932924741693, -0.388467108405254, -0.325053305454397,
  0.045395194457719, -0.593371459992757, 0.352316935904806,
  0.504737258512463, -0.248156473634298, -0.342060514937016,
  0.18283010860248, -0.0794711521873945, 0.302702033433285,
  0.171005564761866, -0.593918825859667, -0.346033985918479,
  0.648803145662075, 0.135601400662304, 0.713393648117024,
  0.176590444222394, 0.0777015385100837, -0.0751572293950023,
  -0.00863611010573502, 0.332316340712688, -0.396381600468317,
  -0.792849631465127, 1.87436966985811, -1.13229479907859,
  -0.240046057197251, -0.371166497387274, -0.406264442651013,
  0.575317114358114, -0.67261691397578, -0.991882786278324,
  -0.129050301957831, 0.194309667752463, 0.283674507827442,
  0.272690613168295, 0.149903179549589, 0.0996772652423999,
  0.083463061127261, 0.108251207777584, 0.410642916412001,
  -0.158816866348957, 0.26880906461702, -0.336924269199918,
  0.0512328404657757, 0.0362724685746034, -0.0731448165300756,
  0.955339762419545, 0.305108456770587, 0.365769885277231,
  0.112952480672082, -0.124058729806058, -1.04620910290549,
  0.349010978150805, -0.0112218549423316, 0.0446401290040203,
  -0.0822668379507977, -0.673973438995484, -0.248275493923031,
  0.599300461194193, 0.3888733576664, 0.155225602366991,
  -0.381678114521454, -0.0943515798031134, 0.272767462470197,
  0.266787470852678, -0.089279258859033, 0.823254821129637,
  -0.464161475796599, -0.471259566908832, -0.284035409001012,
  0.172296128364378, 0.0747712968665784, 0.023163327256444,
  0.055239108176888, -0.27730873318101, 0.734815257867247,
  1.3226054966971, 0.447218634773633, -0.493696566084698,
  -0.150008686930579, -0.0570478084338275, 0.0476384090699624,
  -0.222520552902962, 0.193153281254349, 0.00373244769843405,
  -0.0764502859838587, -0.180188842489548, 0.0375662250147072,
  -0.0201610354051861, 0.0939540897594524, -0.146054480868606,
  -1.08759035086553, -0.578676083600097, 0.795922044109556,
  -0.414413291380027, 0.414190223975614, -1.36156112342065,
  0.225687107294853, 0.169381359108523, -0.161943765171176,
  0.220681859218058, 0.0891683069291329, 0.270994651826449,
  0.465691683840354, 0.518119872554727, -0.248525951427768,
  0.212209719812661, -0.0428753501682076, 0.257452144852828,
  0.205477875725139, 0.0926323581317078, 0.173512833994327,
  0.673847103859123, -0.00457062861531254, 0.17260690523334,
  -0.438921647532022, 0.0844826528545307, -0.173541777088241,
  0.0548425924175375, -0.309583296886564, -0.286765596630369,
  -1.01993275154003, -0.258602477743505, -0.238922685709216,
  0.177732339081788, -0.0261156230798717, -0.162704003581286,
  -0.43219379412686, -0.532586283102987, 0.572638893113759,
  0.238570102092811, 0.558580588948277, -0.0594297125594495,
  0.119201837097721, 0.109728971601297, 0.357265611759065,
  -0.121510488754509, -0.177420139165373, 0.476179279588833,
  -0.543885234637891, -1.00564683322902, 0.151946736106525,
  0.0876480659766223, 0.0835428412369693, -0.189946306132917,
  0.228214281780588, -0.562920583747734, 0.0895589369943568,
  0.505328685823619, -0.336456984119422, -0.118076797485996,
  -0.0624982979683399, -0.00950230173495947, -0.167154452136035,
  -0.673938882617692, 0.34394119056791, 0.0592562047262039,
  -0.239357265787291, 0.652743630280306, 0.17244249239088,
  -0.00415931431770699, -0.449029698836652, 0.0935913626295644,
  0.232271082588992, 0.710165754903856, 0.76974043043327,
  -0.178041665064731, -0.0493960588772525, 0.749376799652261,
  -0.132225038196524, 0.0339991141397525, -0.138350539549074,
  0.124807331983443, -0.258424186370781, -0.13404287489715,
  -0.0629459533278307, -0.0117136657448061, -0.191988319250172,
  -0.0552804915071224, 0.0216411936163243, 0.155340251082966,
  0.154435192577301, -0.475650983932599, -0.237872909489891,
  1.02862201344436, 0.202734439328719, 0.535011702964028,
  -0.146990812538508, -0.327226560150739, 0.250023915656496,
  0.222455312567597, -0.474128138193893, 0.276574523208439,
  -0.2852370497694, -0.506308068796243, -0.0670299641236253,
  -0.0205232175603255, -0.18141209419232, -0.0642572822322036,
  -0.31143913106657, -0.0112745322823956, 0.167133079427386,
  0.181915130773026, -0.602635765864769, -0.545881524495274,
  -0.0216308030922603, 0.0188629560934867, 0.251423879831653,
  0.653128609657551, 0.0629478849670894, 0.333297590151695,
  -0.198049937686654, 0.87877281648551, -0.643343188405701,
  -0.147715773372467, -0.354445905222437, -0.105602168092562,
  0.0442567144641517, -0.682419267000423, -1.07575120295021,
  0.173671056549046, -1.17888450770657, 0.512466965480139,
  0.305081490250596, 0.212103091986366, -0.0586707649680639,
  -0.388781420871126, 0.222546166809004, 1.07517762193601,
  0.925268985287074, -0.414720710549807, -0.0776908147389364,
  0.217071485789988, -0.168757323985504, 0.140610758727301,
  -0.21546447238908, -1.46724425941937, -0.374881689850677,
  0.647752019117852, 1.00520854910999, -1.01734789517651,
  -0.46898590293566, -0.0504786652262511, -0.182704871935315,
  -0.174035574889608, -0.146269900580442, -0.423276567098593,
  -0.546358206909698, 0.15433245719686, 0.28787823180325,
  -0.093440113525012, 0.235993105254384, -0.0339204338279253,
  0.0657611405288588, 0.197451254972995, 0.919741149558016,
  -0.181385028744711, 0.162049876466857, -0.983427008781317,
  -0.0964025522688768, -0.122637147459252, 0.11580717490253,
  0.211502704500486, -0.515664410511978, -1.15036295834799,
  -1.14118076487014, 0.663557022927813, 0.158666344036876,
  -0.450376053309847, -0.172335969050841, -0.0392610365294117,
  -1.19882244255172, -0.195488789861999, -0.288166355971453,
  -0.292934423064576, -0.449411674852618, -0.300232076169726,
  0.105025136810359, -0.0578599458525187, 0.180516366098565,
  0.220023015523402, -0.108002383471825, 0.204264768944278,
  -0.257710481062408, 0.244197113228451, 0.693369774468212,
  -0.0650392297232139, -0.209907683573699, 0.205204711131405,
  -1.73420023203776, 0.733885462203378, 0.13362469131054,
  0.401986402978079, -0.0865756056496294, -0.734919901058754,
  0.295759110556236, 0.0553146832120991, -0.00790075374427771,
  0.268054645148968, -0.252962272938845, 0.536380007483555,
  0.335402415562376, 0.455983818864536, -0.74839176150716,
  0.15383291808201, 0.0986619490301004, 0.205138538890498,
  -0.720010867739358, 0.0163132982386538, -0.0936407932560159,
  -0.621089218021024, 0.509972744668372, -0.418649481598149,
  -0.334469888515089, -0.301549052740708, -0.30225910837971,
  -0.888085079703354, 1.05439381654749, 0.235784473748875,
  -0.637429445246174, -0.368419355595961, -0.585720493864606,
  -0.10276307302283, -0.128608712252482, 0.0582440060390023,
  -0.0143085162260421, 0.307614603824201, 0.468536675647434,
  -0.266042997916635, 0.187936178034787, -0.473472876888982,
  -0.0306735762654407, -0.136062543002837, -0.031412117370624,
  -0.0368330299562993, 1.78165987999934, -0.116511310971268,
  -0.251470139091375, -0.323163910620768, -0.020769327708855,
  -0.0546973577219891, -0.0474509089577824, 0.329793691710631,
  0.0847977075382167, 0.17785507818963, 0.0737711593965529,
  0.834341781618318, 0.769838559776787, -0.524859055632111,
  0.199989370680443, 0.297135078360887, 0.0318278800514649,
  0.315116293293244, 0.554337283060816, 0.238190539516097,
  0.250179006988239, 0.163537760686534, -0.0125637520618844,
  -0.0537998117175399, -0.215337366005561, -0.0516059860110268,
  0.700436682902202, 0.00744632033222245, 0.0279393244705829,
  0.397499248031972, 0.154892080921369, 0.40645513182202,
  0.123497632028426, 0.0122014488165258, 0.121024483234685,
  0.410597477121462, 0.46994752903513, 0.521967253109114,
  0.0504703944271752, -0.754920342743898, 0.0964207226930687,
  0.102504971984811, -0.236133084795529, -0.235416536384787,
  0.254187218642758, 0.420102541914657, -0.167158245339337,
  -0.825996305711818, -1.26861087092039, -0.302839462855569,
  -0.036167495723572, -0.703341191406326, 0.00540834525816589,
  -0.793303186213366, -0.0472207066781423, 0.553523299161916,
  -0.637598477099041, 0.281262900538205, -1.32914951961674,
  0.189320169414496, -0.190518812706725, -0.0432233678646741,
  -0.894706714968379, -0.559750354070958, -0.103738484914558,
  0.460738245462511, -0.346594697116096, 0.0479206159171142,
  0.129306326345626, -0.089243911302499, 0.0119581934711552,
  -0.713217373676302, -1.01024850501196, -0.175213087913461,
  -0.30323536355208, 0.705491689341158, 0.916784618533583,
  -0.0124711048506637, 0.353140369753705, -0.153006211205361,
  0.174001927253248, 0.498945920476948, -0.799178498655451,
  -0.22709656735592, 0.433504296208465, 0.620940037333123,
  0.233314332013937, 0.0935814809066603, 0.262385981559604,
  0.585109129872773, -0.666091561389166, -0.349582021720855,
  0.894513819329093, 0.632064496931137, 0.653074248510619,
  -0.143854014688995, 0.215158132269324, -0.0685703828233301,
  -0.0118877903202885, -0.151436712214121, 0.122044482847441,
  0.115452451257065, 0.210169080685667, -0.28912827169772,
  -0.242354658231993, 0.205830240464313, -0.122655978194848,
  1.04024204968691, 0.665253362828192, 0.759135026110759,
  -0.133048291489758, 0.241035274503402, 1.72264877069e-06,
  -0.149837314644642, -0.179889727036156, -0.175835198491446,
  0.918381040270623, -0.493780964671473, 0.32439158030945,
  -1.01545221951647, 0.0534875198410291, -0.440569555069818,
  -0.0956624788620444, -0.108163170604454, 0.361670887608888,
  0.134630381848682, 0.332615287614696, -0.214432519438502,
  -0.131596879676686, -0.333208439933604, -0.250324308520353,
  0.111486146295008, -0.198595243145086, -0.267659100589294,
  0.231971766484696, -0.0479052057348664, -0.298640435907665,
  0.117390366347726, 0.046804077801938, -0.466355377150121,
  -0.210024025624692, 0.0484216754081308, 0.0984572721747181,
  0.679010766319547, 0.440813874144537, -0.279770069718393,
  0.63207021113297, 0.565902518825172, 0.0102902570469086,
  0.174621747662896, 0.0114013734359081, 0.173143829116808,
  0.276588487265314, 0.0327735163296421, 0.195967632319219,
  -0.559838637155161, -0.106652997757146, 0.238843700737298,
  0.0569306132196164, 0.012810950026766, 0.0382663410118889,
  0.782352676677517, -1.13537809313479, -0.556681075453618,
  0.462339066746695, -0.500939394868922, 1.02067890980863,
  0.0358981868975053, 0.0537197824263473, 0.178250643338022,
  -0.110160249241086, 0.330318529471281, -0.241719175143848,
  0.712557048060339, -1.04270759053015, 1.02408612868395,
  0.0222274207740295, 0.168733491186156, 0.0690143346801109,
  -0.219033102622464, -0.0304221358599985, 0.266347114514435,
  -0.00570296246931685, -0.619143172946276, 1.37336597344578,
  0.147428509079949, -0.228950145791917, 0.129439316490034,
  -0.32375705554806, -0.173459096740565, 0.166387994749522,
  0.298106692000113, -2.2399373357218, 0.299624552987906,
  0.22030343779421, 0.310603574863077, 0.0478391969825307,
  -0.0907085706044047, -0.906283666655288, 0.131337789476489,
  0.326483991520812, 0.881254099171887, -0.107869341126581,
  0.112382955063041, 0.213076584728456, -0.233785423619847,
  0.509170141272205, -0.089428655045853, 1.26841531915043,
  0.0266637192163053, 0.410974261327665, -0.62059005383644,
  0.0712604086502553, 0.0458336983572077, 0.150869186537682,
  0.0625337330536087, 0.0531454168301918, 0.168908069946079,
  0.637171045180442, -0.0647912085765966, 0.381764204168677,
  0.0460969996921838, -0.0839724052296568, 0.0562447664988386,
  -0.471530211406677, -0.928541274171454, 0.857185326574836,
  0.828374437243785, 0.762876144865797, 1.81556134059004,
  -0.0962383856590017, -0.082146245214056, 0.437305123256286,
  -0.0259722464646497, -0.56257186466237, -0.42419393970943,
  -0.3308990015734, 0.0593721593037062, -0.380681107009722,
  -0.218298421818067, -0.00511469068761255, -0.240323387623302,
  0.877507778120805, -0.63450064981966, -0.999510295465824,
  0.0812576357296497, -0.480818661844337, -0.557269393861281,
  0.0509158199405584, -0.30510460459849, 0.0026377519260922,
  0.110071895756987, -0.0716280589696346, -0.407544613242019,
  -0.279433280672918, -0.566895238150737, 0.315482827385276,
  -0.187906202938078, 0.334813725120546, -0.0162925175187457,
  -1.20562459068292, 0.31646220194412, 0.808535906224379,
  0.00211832160065301, 0.595005479377176, 0.170473179932556,
  0.314468596594482, 0.0482749393779111, 0.0581315436041461,
  1.29640801569775, -2.00891692009327, 0.239392840012342,
  -1.33461818112088, 0.810447383940183, -0.520069963629458,
  0.243808428643653, -0.362528480721391, -0.0921798204913966,
  0.254999683994203, -0.242064511498683, -0.443183352792233,
  -0.313105627701536, -0.22728170796948, -0.407864967688811,
  -0.308409376218891, -0.0467349698474233, 0.126293440464987,
  0.233299594781833, -0.267481854876687, 0.0294947507492256,
  -0.0352496986381347, -0.230713424274472, -0.0813802119407066,
  -0.103203095302514, -0.234122340605828, -0.0411502683106342,
  -0.262199637055932, 0.361804700308466, -0.740620852427173,
  0.636695409618706, -0.862203945260383, -0.0450914932572101,
  0.0940406634904442, 0.309092008158187, -0.189782567478971,
  -0.666753604846772, -0.736658159332911, -0.0730436854955585,
  1.17331157951997, -0.229106736078606, -0.618885416428932,
  -0.167654738003424, 0.0638536057538162, 0.0624381395223322,
  -0.290008060863436, -0.794501196804631, -0.199999939998427,
  0.100021729442327, -0.449169467557544, 0.536786485459568,
  -0.0664972551956442, 0.148700706657283, -0.0339493676422312,
  -0.113267454635352, -0.861522961862603, -0.384281565692584,
  0.095813965531897, 0.229888159088123, -0.219811456945668,
  -0.0193244011485532, -0.00950915526831724, -0.259457745804468,
  -0.423563208562541, -0.777845044747505, -0.0923383816290215,
  0.93862426241693, 0.292434328603782, -0.239811494549665,
  0.0573756489904959, -0.0398090201404784, -0.225690481557573,
  -0.703279804276047, 0.516140632693643, 0.401515994120109,
  0.259845502489232, -1.37162855167725, -0.507832379086934,
  -0.0519196220990936, -0.00364634828563412, 0.251466008317225,
  0.59373079730345, 0.206981882478353, 1.27053290884513,
  -0.784299388515554, -0.336398070387103, 0.0764638230385918,
  -0.0168951876452224, -0.166576105912129, -0.228291385440463,
  -0.303666501229496, -0.168657285225513, 0.211969298665448,
  0.207961738061994, -0.0479982545387276, -1.12026920670403,
  -0.608591578765604, 0.155440032278902, -0.0912705720879475,
  -0.895155655156134, -0.310701798740301, -0.845925238079773,
  -0.0611906145057307, 0.11053712785399, 0.0845673409268546,
  0.315482504116772, -0.0207695111914493, 0.236269093412668,
  0.101340916105773, -0.316891153512885, 0.80417405093459,
  0.57533717605836, 0.526371834875922, -0.754694208675693,
  0.0224847409470969, 0.0566191963466978, 0.409973244686318,
  0.248230957000447, -1.17998205693673, 1.84968086838415,
  0.613271755540026, -0.600998724019218, 0.652885953056484,
  0.000935018506684521, 0.00707529099000963, 0.0500536822052285,
  -0.401581606847951, -0.264122265316175, 0.451340668077159,
  -0.279497322415782, 1.04560005282143, 0.104579914236691,
  0.247256173961858, 0.032086385256322, -0.0403650294847613,
  1.18305706350573, -0.413481294988115, 0.30811203864086,
  1.27777742155936, -0.678288146522081, 0.323744439765739,
  0.344077123452326, -0.346021529429123, 0.0778191146850565,
  -0.564947342162814, 0.313465929479075, 0.400093075836688,
  0.630488174397964, -1.12968472441505, 0.596010993823688,
  -0.325207552400236, -0.19771617305145, 0.103500754358472,
  -0.293093555607086, -0.660096438925857, -0.332105423647642,
  -0.223988732045849, 0.201817359497599, 0.251637676072312,
  -0.210455814155953, 0.239600175204037, -0.0651207430477812,
  0.373186643302469, 0.200169738753196, -0.083349315236508,
  -0.294833737824635, 0.318460398552108, -0.387480637362929,
  -0.214783293612065, -0.0840994234127382, -0.0981268069976287,
  0.540527161055998, 0.022904405138292, -0.255378572724474,
  -0.197705993334278, -0.0512506874059647, -0.540884628815511,
  0.166512294575122, 0.0554734844132567, 0.164848819317236,
  -0.0678145392693225, -0.465898339994158, -0.131493033699191,
  0.938942353377471, -0.418238367675548, 0.148672915566515,
  -0.196402187176935, -0.195367974526426, -0.0193513714341956,
  0.164881444107007, 0.30447968713302, 0.106507813051214,
  0.26886304455404, -0.288620950027129, 0.0208552247210121,
  0.0116208945607255, -0.092318591218325, 0.0186574842856359,
  -0.292244405780905, 0.222116654394776, -0.042161251776968,
  0.076857425637727, -0.117050183225184, 0.121996391667862,
  0.0211089866708939, 0.339108982132363, -0.26492999461197,
  -0.47668961965632, 0.177369892426964, -0.332150068620268,
  0.497268742199388, 0.509357867540056, -0.143775104091674,
  0.023908501791824, -0.130143292597557, -0.125526803924789,
  0.751068331716108, -0.223780720292787, 0.525616372367607,
  1.31635412859905, -0.268630937334943, 1.05626747412668,
  -0.327497314770788, 0.443886991083927, 0.0177831083914886,
  0.227821808206765, -0.14103517659373, 0.335877578500005,
  1.01076106043187, 1.16531988013291, -0.245515913771667,
  -0.126248473741381, -0.149037317491679, 0.200807567576062,
  0.030336927376822, 0.288631615236924, -0.197790062717797,
  0.36231676380893, -0.157060949980036, 0.687653321461091,
  0.012187694719254, -0.193667472788079, -0.09802397964628,
  0.0104279584925375, -0.302372620119059, 0.0201637558277982,
  0.431415672626506, 0.505356719536073, -0.334792171844074,
  -0.376793229453347, 0.039126313848382, -0.109560766548576,
  -0.642928405671846, 0.155728277023262, -0.394418523693442,
  0.194609908769986, 0.438605617974497, -0.472273056109768,
  -0.0494053411564917, -0.156985668988134, -0.0391959393099638,
  -0.65192244921666, -0.1797970428636, 0.382352445321882,
  0.578052586592273, -0.297341654060186, -0.563418994341217,
  0.0691743219060117, 0.114611369343174, -0.388218855783752,
  -0.215813366299306, 0.0372264170483959, -0.404400095316503,
  0.133261227133856, -0.136892148909783, -0.475534299931503,
  0.0884102990177495, 0.0508221423852722, -0.0655822403823625,
  0.267106842933582, -0.360728221515617, 0.740215873322217,
  0.116310650783663, 0.600514754879824, -1.28731678031759,
  0.00209656772338533, 0.044310480019757, 0.0798613596417598,
  0.597224946537874, 0.329687262816994, 0.606398463370479,
  -0.390753786131069, 0.253443444178947, 0.430060293801693,
  0.292546777376105, -0.162683085642328, -0.298579796412067,
  0.542688863026254, -0.509611561363722, 0.347660188820262,
  0.424971565204495, -0.235368409175711, -0.295105703181304,
  0.136612056988308, 0.209518729480615, -0.242204825692082,
  0.336751838402349, -0.196061099290941, -0.102762568911278,
  -0.0933368582674942, 0.116167814745395, -0.180515473887889,
  -0.160723636884311, -0.0807513276153584, 0.111470463660611,
  0.178531003376746, -0.263879521988165, -0.228136272541203,
  -0.825012807647516, 0.388217171997639, 0.802353006127347,
  0.277434400500989, 0.213790265354674, -0.170522938367404,
  -0.118401298062719, 0.166025216271328, 0.476280217202884,
  -0.292159785458249, 0.101347884250837, 0.440038656610285,
  0.217978279451348, -0.243030929399753, 0.110466366197492,
  0.260781387894181, 0.119206507818176, -0.370383899430993,
  0.765965461218741, -0.94723962376398, -0.207672107619091,
  -0.255853563172774, 0.0112474260724115, 0.0358494318914869,
  0.0126221222043473, 0.320578851229126, -0.209279709433274,
  -0.850536157084454, -0.218685999657088, 2.06441319363544,
  0.0581078085592218, 0.21654121779202, 0.14999133620141,
  -0.435821090432815, 0.273821733599542, -0.451482485261147,
  0.288840623893277, 0.528360385041737, -0.0376893358201596,
  -0.192651790702306, 0.510341300103034, 0.0921636109173079,
  0.101063556190114, 0.466250884055339, 0.259189904919117,
  -0.451082538123625, 0.467529581824557, 0.315429134822411,
  0.0307373662892918, -0.0974157940819672, -0.195356839810604,
  0.478454122347757, -0.481941457586592, -0.138511387235107,
  0.255512755943431, 0.227295678504522, 0.661570597917944,
  -0.163326327303334, -0.255342408405753, -0.0378076714616273,
  -0.223351112940492, -1.2061156911942, 0.0164228243373308,
  -0.993226398113614, 0.705502503621659, 0.583954831926191,
  -0.047131895944726, -0.284701017516458, 0.0120442671877007,
  -0.0284319521093218, -0.758333278131147, 0.135463877513586,
  0.360041838864735, -0.759835777548602, 0.0265750848519362,
  0.214042354329536, -0.139358858988957, 0.33499148732382,
  -0.40955287118103, -0.730002877740021, -0.307106735307693,
  -0.359045293480376, 0.463441053755317, 0.785783210393286,
  -0.269394967711897, -0.00121143077904325, -0.482159408542053,
  -0.0600096178858049, -1.03021796336695, -0.74451339088441,
  -0.948258936294937, 0.346583235476973, -0.433276725970432,
  0.0816324090789821, 0.125287410699396, 0.0798307370394922,
  0.20262003237656, -0.224799164737478, -0.0221888497793247,
  -0.193594002862621, 0.450434673363703, -0.403570538699052,
  -0.166336291627812, 0.0866190164087418, 0.277926720111462,
  1.03559677725618, 0.724303376307088, -0.124190944970136,
  -0.830903804241739, -0.740191667606211, 0.617750724125057,
  -0.0499631202717255, 0.144910227580966, -0.0480947973671049,
  -0.430156366075413, 0.934226641997182, 0.672832379020635,
  -0.633510327841067, -0.499079151674412, 0.270353927893189,
  -0.174359377008032, -0.286283270787299, -0.0619058795767706,
  0.0828442897264522, 0.527023435861187, -0.111486214281408,
  -0.775631296094406, -0.840654997323189, 1.00266301652195,
  0.212162301552224, -0.251934892146406, -0.0253081700149028,
  0.957654661299891, 0.117603078577674, 0.925570795943348,
  -0.116798630875436, -0.403485372735502, -0.180183034311058,
  -0.0300772833868071, -0.215666170394519, 0.0657340352155201,
  0.523514449936676, 0.0388771009449598, 0.215692542443473,
  0.0581141525640511, 0.0313034170011113, 0.0601638863980312,
  0.260947498972336, 0.175827447845638, 0.00145502784338618,
  0.394163641608694, 0.0734111953331292, 0.0603698752836882,
  0.401036871821251, 0.472097769191558, -0.244622750773965,
  0.150965451902855, -0.204221487437509, 0.0853469173527346,
  0.254378280402159, -0.307743016487218, 0.213989808543307,
  -1.3256072808345, -0.881149730691815, -0.975609684739828,
  0.14946508756845, 0.214080813740026, 0.125071304143361,
  -0.12629251852059, 0.123277743299782, -0.563329086177585,
  0.0658966222775174, 0.745682365997224, -0.11069608321231,
  0.374514820555116, -0.155637891139439, 0.30512196279904,
  0.268412841767102, -0.541696536469414, -1.27608278629139,
  0.0252552834315531, 0.659509099648122, 1.26389673288762,
  -0.26678659631126, 0.218215486853975, -0.0314421911580887,
  0.152123888147941, -1.03792173325059, 0.273903268697355,
  -0.24659339818282, 1.00339110587492, -0.183119981617482,
  -0.136165774566811, 0.0477389495416002, 0.354437276204049,
  -0.449935558967739, 0.507814459289193, 0.498742767772381,
  -1.14952823718063, -0.603360611415992, 0.62527845631162,
  0.106378873537953, 0.0262284934231398, -0.112929563830579,
  -0.272904853167294, -0.155344289958113, 1.81870347216707,
  0.156679126795912, -0.295803726052628, 0.699121905000203,
  0.23029247106236, 0.0153897566598323, 0.02332786139659,
  -0.238101260642007, -0.227107804768789, 0.0988624077359397,
  0.104969681879671, 0.252213236363577, -0.299774784825046,
  -0.100577708039137, -0.239454545271328, -0.3511659503874,
  0.225612540558428, 0.985241541602814, -0.952689669562297,
  0.212558111469693, -0.893021292261741, -0.585729807392702,
  -0.334143047792353, 0.00198548616380148, -0.202416841687917,
  0.925215389320549, 0.167250410641958, 0.356668782875545,
  0.0288420927666609, -0.0981661442013857, -0.237486230171152,
  -0.0283917306409919, 0.141579374344261, -0.00262174872932341,
  -0.071694824536229, 0.164135829162007, 0.736888386413375,
  0.186028500443998, 0.0784490738351664, 0.616604829805622,
  -0.0277011930248438, -0.266892638516401, -0.0149615507402762,
  -0.282256864721236, -0.404051665993076, -0.849062396854254,
  0.611954374486427, -0.414962348797283, 0.680026223209408,
  -0.244727823351837, 0.0447515314334728, -0.206394671133311,
  0.0780508441615234, 0.0287653404072076, 0.647806479503341,
  -0.374348129510825, 0.536753519477371, 0.688100925931323,
  0.215994108658542, -0.17503908430497, -0.293906103244192,
  0.20914205729631, -0.541541463272316, -1.12458095129547,
  0.195217381706786, -0.419490922016281, -0.780832036880052,
  0.190287432630335, 0.105242878470342, 0.162673184055686,
  -0.510215524160507, 0.0476028313810591, -0.321011834013036,
  0.349367126342142, -0.684307205393608, 0.528671771497834,
  -0.0860504414560772, -0.122062578838156, 0.318923874963348,
  -0.672805674569334, -1.11811092499164, -0.691038723607512,
  -0.214541458783806, -0.231241493575798, -0.853105618314957,
  0.189497416647639, -0.084489512101431, 0.107839451938501,
  0.81219454473086, 0.114756208151743, 0.509668286454313,
  -0.0864222071484341, -0.240469970236505, -1.05443053151225,
  -0.0356887231240274, 0.00901632043359718, 0.15806939134072,
  -0.197144163734535, -0.33612311719493, -0.161530665826825,
  -0.443963302750047, 0.276661212226422, -0.380886102079002,
  -0.405216393319399, 0.343336567911506, -0.0314958541084642,
  -0.788127440505554, 1.32388450203935, 0.0483299180835698,
  -0.367907192064245, 0.0436021247531413, 0.490519740594177,
  0.271684765563734, -0.0415262559050757, -0.119229468533045,
  -0.357120920403137, -0.211438816091911, -0.232574610906385,
  0.519710070021466, 0.0831045883416086, -0.40449458966511,
  -0.0775872725862851, 0.0211768047340068, 0.0477652319945192,
  -0.42717199967403, -0.235041850221706, 0.186456093309766,
  -0.00758034108300306, 0.171087101758743, -0.947175078184485,
  0.126957229265181, -0.0115062572296736, 0.324314936214408,
  0.212252601717993, 0.0268702250242775, -0.235650341911832,
  0.135184015106446, -0.0552999076660499, 1.12906198435448,
  -0.124865232451773, 0.0159904531005839, -0.162575114096937,
  -0.403124729527502, 0.877041713052347, -0.695991790292825,
  0.31411543932363, -1.3047239745879, 0.652742784033591,
  -0.191151974966988, -0.171577836929953, -0.0747205734507797,
  0.582495968233043, -0.263388227221216, -0.431378392016922,
  -0.415448408943933, 0.18804086049976, -0.579092049804233,
  0.193068618623397, 0.0397558573756717, 0.050045994899123,
  0.195796409975254, -0.244160937748033, -0.658545056487517,
  0.215501169434917, -0.186754330196084, -0.340903013319281,
  0.426621989754263, 0.0790322615412185, 0.0904919584896798,
  -0.769344333461963, 0.181148298018301, 0.23216672392847,
  0.246676228890354, 0.539441317520061, 0.123637276409115,
  0.112020869037792, 0.205506264396656, 0.0453531832858616,
  -0.333950290167439, 0.0901436044847694, 0.211223604955023,
  -0.66534611018078, -0.00655916320350751, -0.214988506277981,
  -0.00258564273676387, -0.25395091623441, -0.0651303668657735,
  0.330925122138683, -0.478649924990973, 0.266143964630676,
  -0.224429350274322, 0.324248759070218, -0.313550442810772,
  -0.283699031868329, -0.183845439477192, -0.0202794119155198,
  -0.42959759704301, -1.13227038812197, -0.441627831194222,
  0.0758824326365819, 0.252113975292708, 0.386956284170888,
  0.0792682854056682, -0.174941179543674, 0.188077814301803,
  0.102109856181241, -0.154606760470825, -0.0324100037860309,
  -0.0375971828370798, -0.223892355535361, -0.639748633009499,
  0.11521996398232, -0.444025575773755, 0.0569865012429926,
  0.450792206260931, -0.832505761410813, -0.260141255183714,
  0.912200296178486, -0.70479959879869, -0.796034363403832,
  0.215504239417828, 0.0101019833747244, -0.0625187048934426,
  0.892391512021768, -0.541093062767475, 0.485041195361636,
  -0.542152116901785, 0.450515817235422, 0.955160957890025,
  0.0471624330051861, 0.254857961176274, 0.183897700228555,
  0.904130261622563, -0.635254559624013, -0.496897453959245,
  0.371690088539729, -0.689918183214352, 0.561502941351985,
  0.114559469260615, -0.12061031369704, 0.222619010303591,
  0.409817729052443, -0.423965087409404, -0.0682788773349166,
  0.307472962374921, -0.0213727146497229, 0.0945842852698404,
  0.296779717046999, 0.00772371049874759, 0.0220674327618596,
  0.790006822390794, 0.0515516833193047, -0.156715125121881,
  -0.309757222291325, 0.0762206840561225, 0.892282663629755,
  0.0184784489363696, -0.290666381271613, 0.0636853061553158,
  -0.671763302912732, -0.19080018491236, -0.217260395627206,
  -0.527481833645548, -0.149258384616436, 1.20599845392024,
  -0.0134293349841187, 0.0644302297610567, 0.106544312631475,
  0.676825754599756, 0.35972396671078, 0.0865689864637216,
  0.315890217208936, -1.60747922361851, 1.58301158767755,
  -0.0112314958242916, 0.264331783131261, 0.531426712142776,
  -0.639533084003201, -1.2026842122467, 0.301107879360298,
  -1.20571280947046, 0.523827909385833, -0.633927868569543,
  -0.238911112589915, -0.0957122310578023, 0.0992237349075828,
  0.7583422584048, -0.413245111163983, 0.282169246413397,
  0.187954065676474, -0.378770470696185, 0.184862497546211,
  -0.051689437624272, -0.0474568753626424, -0.152603312017219,
  -0.753218780189194, 1.13024139976063, -0.354501914562605,
  0.30849935670834, -0.327248888955928, -0.195856961595942,
  -0.172665836416595, -0.302019884897088, -0.0610128299588322,
  -0.197832335230087, -0.275735977256222, 0.0327907186141723,
  0.0732386787073691, 0.0669531850060115, 0.251351728894157,
  0.232175189330325, 0.622444303433632, 0.114492190289042,
  0.381466637890674, 0.63470706502527, -0.0592036829467147,
  0.029631059771667, 0.552286990329221, 0.514034167229052,
  0.0251797486335382, 0.0695596536248735, -0.0177474892429768,
  -0.0629100046794976, -0.102687457236946, 0.270281306664286,
  -0.144737648182441, -0.543615124891365, 0.159361822643806,
  -0.158575334944764, 0.0370900557017594, 0.0969598515335886,
  0.32309526451178, -0.0143802446569884, 0.309201812944456,
  -0.158592924639043, 0.0115598003286322, 0.115297722107069,
  0.012392307606522, 0.322354875965393, 0.19503571715092,
  -0.0346008769092888, 0.949524926784433, 0.0825869321378213,
  0.531992738439155, -0.230712255516604, 0.00174194006189225,
  -0.0278841618613188, 0.0444803970263118, 0.167409788659322,
  0.172066945157166, 0.307782456429489, -0.0149566857668856,
  1.10936335702296, -0.559129021054405, -0.318091430607124,
  -0.136668654385958, 0.0973283479183581, -0.0578681366954763,
  -0.251276599773947, -0.963008690877286, -0.247652635882225,
  0.348101445660525, -0.0213843824764647, -0.614328726692037,
  -0.095931903061576, 0.386293410960654, -0.00594371592196152,
  0.393843552887247, 0.706282444255402, 0.491146364987031,
  0.00472197919627925, 0.454458330522658, -0.0893737202741318,
  -0.150938128071746, -0.0349490226591884, -0.0639840003763608,
  -0.437930471977602, -0.304257392915743, 0.347640995155652,
  -0.124753585160887, 0.48201509577197, -0.00631010839488878,
  0.0381632029891461, 0.0867099145368656, 0.192122551653241,
  -0.276940764668586, 1.29785506673055, 1.02240448491423,
  1.34367767646621, -0.39786921213819, 0.0603222848969222,
  0.186472648482914, -0.0293728734239046, 0.142072191709634,
  0.660675027014921, -0.269619101983582, -0.0306558548325262,
  0.124873827975826, 0.339734966638062, 0.157990945573301,
  0.136180935995707, 0.0124024915526498, 0.110943234012334,
  0.473483908724695, 0.121698161332788, -0.320152468429535,
  -0.0183021582422652, -0.305223944425335, -0.0456368048824794,
  -0.152049073721807, 0.137019570427255, 0.139737783394691,
  -0.0948245554505168, -0.72054219083962, 0.0763830568932191,
  -0.111892112243522, 0.0927657048714364, 0.213811157287287,
  -0.0877923270635791, 0.3916623676173, 0.0410105029934351,
  0.328407191743685, -0.434802587903557, -0.416848190915508,
  -0.208092717661381, 0.711667677660823, 0.325393407939196,
  -0.169501351619282, 0.248695498176488, 0.211927842784388,
  -0.549380072471379, -0.337748946297218, -0.43507268722407,
  0.360758083320631, 0.376602008381615, 0.00757839812707899,
  0.210424445271918, 0.27610432162756, 0.310265082526302,
  0.284908545156312, 0.135381143129556, 0.514397429228191,
  0.608538917678402, 0.202493023788324, 0.386405219268409,
  0.222939640207141, -0.250914066500017, 0.0750522333331398,
  -0.042128061129725, 0.358082531602095, 0.068473873993146,
  0.41408556185288, -0.735820367443738, 0.14743265059335,
  -0.111645946160594, -0.0826808835608933, -0.113777454632088,
  -0.963153286250652, -0.355974849719056, 0.533887990058212,
  -1.02458812085299, 0.978243031600147, -0.542469180703935,
  -0.0862728934033769, 0.0855484642625026, -0.430045604158237,
  -0.141857108938518, 0.597985649467121, -0.749759548452144,
  -0.572280268720761, -0.13860700047945, -0.365185483711128,
  -0.109307892726463, -0.370472467477678, -0.417254778250838,
  -0.990951792810916, 0.149635350504475, 0.222665115505975,
  0.702682273858017, 0.308610255382966, -0.469042458985533,
  0.0160447462946805, 0.170753381238013, 0.0159990303771844,
  -0.216979428166018, 0.064801141000789, 1.17648417177507,
  0.252889294348412, 0.817017081993839, -0.254420753540905,
  0.070862736730298, 0.206275791543329, 0.0383905306056669,
  0.246211328007176, 0.562421234702544, -0.105680126728833,
  -0.623631593317889, 0.217702063448444, 0.463328500905331,
  -0.0449385543290162, -0.173157429881723, 0.345522739744764,
  -0.132713853558638, 0.18186806415467, 0.13315708106165,
  -0.1494067558342, -0.0421408047312764, 0.351421551279827,
  0.466423993167033, 0.372561971259693, 0.0298177258440161,
  0.0112421617375297, -0.299957436621121, -0.54057400030895,
  1.25268414723476, 0.629195627627385, -0.374361114630515,
  0.246125798165503, 0.030591156243532, 0.19950329128137,
  -0.870585999165635, 0.174102470097675, -0.527009838793925,
  0.524926537605275, -0.17786827522804, -0.36700967987041,
  -0.281348883487128, -0.0197909416404437, -0.17267191484431,
  -0.464268558620089, 0.329876078217537, -0.333424312940268,
  -1.2175698881174, 1.09358652768681, 0.155043400158104,
  0.094975591859329, 0.0718377110518635, -0.0927767308783887,
  0.718161927519135, -0.418131834297422, 0.828903732858027,
  -1.05153255544725, -0.283369132062939, -0.141463509021417,
  0.232656102259663, -0.030292899925494, 0.0872143911662923,
  0.189261852189056, 0.217604908966087, -0.0485664918997031,
  -0.67390932763997, 0.873669867108318, 0.491868706879787,
  0.206442055882305, 0.303285761370919, -0.0216146783598573,
  0.821781257416956, -0.318854801244627, 0.186537765824216,
  0.570310411986702, 0.277750889493171, -0.405184865612823,
  -0.132851056774145, -0.405166210293149, 0.00387718906225913,
  0.693359993824876, -0.0977479473899703, 0.42493030489863,
  -0.992205544713935, 0.271142359368032, 0.205198150846468,
  0.0468670422179367, -0.39306589873488, 0.28948681288427,
  0.3140738523763, -0.614126899022709, -0.0731411756458765,
  -0.466980544934763, -0.735429802724173, -0.0919821732270468,
  0.0594755034094608, 0.180363530816255, -0.269894172783691,
  -0.676559047329804, 0.344496040353256, -0.0278938740787474,
  0.200818273109656, 0.379397589401688, 0.796035774305147,
  -0.175217956728077, -0.135550673129393, -0.505386382813248,
  -0.443303567053788, 0.101834609521099, -0.166978483992206,
  -0.0997134416743686, -0.603220504077284, -0.444430189226229,
  -0.161897742570643, -0.118225011904816, -0.4841767375853,
  -0.178080125720799, 0.0474832825860669, -0.556091965618411,
  -0.248265013489931, -0.108624543818544, -0.628934857551101,
  0.0542785747343971, 0.204756500131403, -0.00447379372621153,
  0.15022054645423, -0.900532696010064, -0.385073940916515,
  1.16281480214277, 0.800100505531611, -0.489308228136979,
  0.110981002818879, 0.645041812262336, -0.0538714558346814,
  0.640794469308954, -0.153051508332208, 0.581124991439229,
  0.764613950966779, -0.342883456797076, 0.750301963643306,
  0.2745177071159, 0.096536490131226, -0.106843799756382,
  0.518558790793204, 0.397558768322545, 0.238489748074209,
  -0.182174235613599, 0.138273340119119, 0.61759451512392,
  0.137660284031939, -0.0809331529562687, 0.374652454629687,
  1.33548033274653, -0.155782206279228, 0.897276664439265,
  -0.357308289718746, 0.991137785818967, 0.347008322743916,
  0.279137056078017, -0.119430827459015, -0.101413295300216,
  -0.220786604681475, 0.50511519463801, -0.705662383231078,
  -0.211630768147595, -0.239638993673755, 0.671532965695712,
  -0.172498965663751, 0.229926134726217, 0.113846601301108,
  0.166274195170691, -0.0802031144684197, -0.00380597742335401,
  -0.45926079337403, 0.261787085216434, -0.330630255892637,
  0.141760644991891, 0.0472567397404635, 0.143314998915781,
  -0.987076647687189, 0.137112194911269, -0.482640570802505,
  -1.29531795594916, 0.272835098734607, -0.852813135278139,
  -0.141210039801325, -0.114808493047296, -0.295034076658736,
  -0.296812749080041, -0.296935804512328, -0.0412292494177283,
  -0.14215793211682, -0.244440466589097, 0.630473881508389,
  0.110110398077762, -0.255435862941066, -0.260542321545367,
  0.0447491576778848, -0.166287870772296, -0.16157381273429,
  -0.160880534931618, 0.198316509916188, 0.272955881888422,
  0.107173694184418, -0.2261671529339, -0.176185046946451,
  -0.563926061064697, 0.541161723764252, 0.267909546358178,
  -0.468403822825179, -1.35187559230567, -0.167431008303415,
  -0.203958659554518, -0.133983797625175, -0.0868217038156745,
  -0.976387541028674, -0.447913450196387, 0.321224231062874,
  -0.138944829391366, 0.460622269682272, 0.050682949978238,
  -0.211609430617368, 0.0209197775928191, -0.12208100421189,
  -0.0245321566819056, -0.44129113896406, 0.538073624000505,
  0.215408523564366, 0.493597338570549, -0.505790126922329,
  0.116794676732554, -0.250629713798606, 0.289912518885218,
  0.229206345379559, -0.426551697462913, 0.945804846005416,
  0.0114033791779484, 0.356950362321625, 0.222451986538414,
  0.0269287511823683, -0.526667770971714, 0.106854647792092,
  0.0966244423711384, 0.120725473689676, -0.248035904173432,
  -0.67409205946802, -0.814167166934187, -0.182342980217234,
  -0.332333472889784, -0.11556267557288, 0.157104660063765,
  -0.770223368308234, -0.123396397332045, -0.970394885347446,
  -0.100998794729985, -0.101811806920573, -0.114246946029236,
  0.330819470850731, -0.107761691256032, 0.0971947877257003,
  -1.42477818783873, 0.43756768108801, -0.154119542813987,
  0.522158397336587, -0.0819826566448517, -0.0784714924668042,
  -0.0546579240087347, -0.28973427782868, -0.0495688773174811,
  -0.788740081257404, 0.596312773394195, -0.022278567306651,
  -0.107482487114545, -0.218378917274273, 0.56546982928509,
  -0.0823877668552337, -0.260026161593042, -0.1664519926581,
  -0.073913379353063, 0.114852541510438, -0.466273539529229,
  -0.17620117457795, -0.347567436879627, 0.0345027230913329,
  0.190054075444466, -0.0201711354487517, 0.143777099564539,
  -0.29197969995513, -0.0422089381536981, 0.693226602462812,
  0.146608755861787, -1.14761836161346, -0.255828370409306,
  0.0905945657144199, -0.0505335786449993, 0.139702478220963,
  -0.148916204755044, 0.329683539484336, -0.311603160636355,
  0.492257566691267, 0.442650373991315, 0.0682384351689041,
  -0.152904019504485, 0.0486290759973157, 0.10359264141367,
  -0.149613302648574, -0.163111214947728, -0.380000437403533,
  0.0354786936733613, 0.570801630634428, 0.00515146943635459,
  -0.0793383063337255, -0.0437643934147034, -0.0337841097329377,
  -0.716119612674622, -0.249770266465261, 0.219283591030426,
  -0.252039895801314, 0.0216487720122812, -0.129220752689988,
  0.0508460985662151, -0.160990391113533, 0.339964172466099,
  0.196809706717371, -0.761965088112882, 0.728382048829525,
  -0.46187105914011, 0.304687241118567, 0.881442301502198,
  -0.193735019509733, 0.05270555549914, -0.34533642138213,
  -0.0385655708632588, 0.279065062323568, -0.473283267447322,
  0.107991894114106, -0.604120300361828, 0.372306513481879,
  -0.0127940176448727, 0.0701160288716358, 0.145982368564765,
  -0.289281859034458, 0.496549991213806, -0.827012718046317,
  -0.00396698433869647, 0.108437817445892, -0.639234671058427,
  -0.0410292893841894, 0.133494672189217, -0.143232633504926,
  0.378743263605155, -0.103704252674579, 0.0763722235748272,
  0.111340117600345, 0.815330126422657, -0.217463403257564,
  0.129518329987526, 0.0304967412094532, 0.160099634197889,
  1.16765900922596, -0.13018160911601, 0.960268304957502,
  0.640919619389948, -0.00667302850695064, 0.711232378644978,
  -0.135326037476627, 0.027182031471226, 0.252350916387476,
  -0.0589599898868063, -0.0702467880293295, -0.25717134523183,
  -0.781687658514184, 0.923268225085457, 0.279333554074316,
  0.0820268961883232, 0.183186528875672, 0.368287072388341,
  0.0637681262414427, 0.13663376092789, 0.360453694695817,
  0.829441766838859, 1.02297612295818, 0.686663251178346,
  0.0622222525721567, -0.287957189685792, 0.518636093752762,
  0.0280912024360248, -0.399870908520112, 0.602279428295556,
  -0.668386071258063, -0.285447324379064, -0.190320657829412,
  0.0184202344315975, -0.0700257729452061, -0.000112484677223305,
  -0.941383319205372, -0.198426559489727, 0.0983153826567499,
  0.605967269785977, 0.109436016319037, 0.727560810856677,
  -0.0889296870385841, -0.235833629322253, -0.257590650067036,
  0.290946355634478, -0.365770018289147, -0.210412545520238,
  -1.13802622350027, 0.648085104753017, -0.509687368994277,
  -0.296018715270398, -0.480899742908034, 0.125965096375548,
  0.871598731564828, -0.76886955395567, -0.407294057990153,
  0.544147296607788, -0.705823416204937, -0.122615236101991,
  0.158027403206704, -0.0769596475588582, 0.03319239366866,
  -0.271512119725295, 0.123237461208075, 0.451268338205862,
  0.27692769379237, 0.480880554079078, -0.333147196121149,
  0.0550712816024573, 0.13193234845827, 0.218236333995821,
  1.2405880247643, 0.56662119715447, -0.719574067617486,
  1.52619138313232, 0.46602153261274, 1.16700480236931,
  0.156193838476189, -0.0998377327538532, -0.0756668305367104,
  1.25250178271167, -0.253324326986414, -0.243309002442658,
  0.348181536212408, 0.135397973624922, -0.108558420540475,
  -0.194839467682423, 0.144253181319725, -0.0572984833319022,
  -0.725769120664025, 0.793455029444019, -0.504405835765448,
  -0.483601413804576, -0.822029873621317, -0.412228033679853,
  -0.186328855042585, 0.0557956420701837, 0.276178132826577,
  -0.125707821149953, 0.638340250878756, -0.80497295746457,
  -0.0286242113372248, 0.324369026242305, 0.23951886893431,
  0.0183365683789515, 0.127995292034859, 0.0807111909783802,
  0.274604144243184, 0.318133859542158, -0.0144138821341154,
  0.982968714756973, 0.565405395027025, -0.151302186711913,
  0.250835778040351, -0.177463912658549, -0.327153939878554,
  1.35918632860163, 0.135497668122139, 0.11850874803038,
  0.233837924681918, 0.775815624462744, 1.10274917007743,
  -0.00820441196548341, -0.288484745807701, -0.146910781859925,
  -0.862298005551832, -0.310138923955208, -0.0850838356089849,
  0.136917189954921, -0.133856784169413, -0.952040334985586,
  -0.0939326171731317, 0.248466680113037, 0.134948532105412,
  -0.594495896699788, 0.381203305567411, 0.341193472610892,
  1.13188159196069, 0.216450998293867, -0.341045045997629,
  0.0373403208559258, -0.126178653571637, -0.183876257853718,
  0.115608925599888, -0.241472660636493, -0.0940463314738684,
  0.119962060083791, -0.0623868936078647, -0.339566927776701,
  0.0723324302094233, 0.153689054675887, 0.307804097952989,
  -0.170874049156007, 0.470600163706648, -0.277280538506223,
  0.111254730937851, 0.0925056686497602, 0.793955432549397,
  0.210027873089248, -0.39322184748754, -0.273355040078613,
  -0.518793164383101, 0.291295597822324, -0.364073523645551,
  0.0624850067740723, -0.444907908164452, -0.358640489467583,
  0.201018970544481, 0.0789688568945751, 0.275545188063168,
  0.381645020176699, -0.0831617595718616, 0.220642712449784,
  0.210876703921602, 0.33346037281216, 0.281225225398334,
  0.442073472399704, 0.0785002659399599, -0.0757419259389881,
  -0.506906884669634, 0.540377456632187, 0.479162865091189,
  0.204336290835651, -0.934964966482531, -0.412875769714302,
  0.19995683140608, -0.0130999736593982, 0.00923557571573659,
  -0.369107303235032, -0.519387805969448, -0.733862599179278,
  0.471691378252493, 0.762828802214941, -0.00847517725270565,
  -0.112559470202644, -0.0237668943277113, -0.176429148716064,
  -1.03278395358653, -0.4572162156811, 0.291557904551875,
  0.706180219635704, -0.140153891425007, 0.0933456322216639,
  0.261550015133334, -0.0843291422247111, 0.151646936068393,
  -0.181707496474754, -0.509019339893857, 0.646664478086896,
  0.263070267775475, 0.575887104089423, 0.709897336102018,
  0.153897771976871, -0.151685737837513, -0.0161089533291766,
  -0.440586813982398, -0.181968207039675, 0.533586960328526,
  -0.0837308014351234, 0.0575884123173852, -0.752213409787462,
  0.0449741094814396, 0.191378400379035, 0.0756116741140834,
  0.0939592628811243, 0.192068840557125, 0.13024997104607,
  1.1912432565162, 0.17696630300209, 0.629896388069069,
  0.212029105817981, 0.0798533816526385, -0.175134271570997,
  -0.29313834252326, 0.345084108386483, -0.777369140851709,
  0.519448704846839, 0.547658332606948, 0.285317960516341,
  0.128248441719849, -0.0709803628880704, -0.349636557669289,
  0.534264120378822, 0.685791911389714, -0.149451749142283,
  0.616603953829397, 0.801220004913707, -0.134855975458083,
  -0.00192443982544314, 0.423692680463103, -0.181747278348283,
  0.408959654231565, 0.537521050918616, -0.311253039683782,
  -0.405619319018549, 0.359501906590826, -0.0748190552815039,
  0.0794317551932943, -0.0698785926436142, 0.0648046323884292,
  1.35737395400523, 1.49261902308903, 0.618108232188722,
  -0.531284546193636, 0.222827099185016, 0.305705143495713,
  -0.0622350595603815, 0.000362936825187223, -0.0130126184789419,
  0.312761317828721, 0.555790786209624, 0.0892705424221774,
  -0.397886219291332, 0.699447619517914, 0.263772236932071,
  -0.0153603271506102, -0.0269284420718756, -0.118760706000943,
  0.768953531492292, 0.459919780234796, -1.62494434161953,
  -0.401772346227287, -0.775895715922214, -0.150565195645547,
  -0.0584059950030846, -0.119995309769758, 0.0329416174159453,
  0.481977091905043, -1.70946531318276, -0.122598038053014,
  -0.356500974467804, 0.939124267304529, 0.361380613443273,
  -0.0636576769426307, 0.224496756970772, 0.130157145411334,
  -0.118996380985726, -0.177925704001768, 0.934386725425723,
  0.142316841441433, 0.691725981804761, -0.793246170819889,
  -0.0569036821332324, 0.039640877609612, -0.211244995098109,
  -0.883899160604465, 0.664745439204415, -0.558186804981762,
  -0.599464299032853, -0.11401430747745, -0.996903069681871,
  0.439635346583665, 0.195803569390291, 0.16338257684672,
  0.468562728155488, 0.151102526496971, 0.566919025522049,
  0.132427406810115, 0.298504104175928, -0.0557864030339223,
  0.0730854550011726, -0.00318334633034929, 0.19449134154126,
  -0.445380952659882, -0.689810356712232, 0.843647881115139,
  -0.0429464026382668, -0.153072199962979, 0.0385422592317342,
  0.162503027595689, 0.00161914726677998, 0.0349940518576903,
  -0.690080773944346, 1.04545537505361, -0.204232519249514,
  -0.81588581867177, 0.252773460703556, -0.550848012523844,
  -0.383714527577509, 0.0706906485384253, 0.110676534293005,
  -0.678377157158646, -0.564447091978008, -0.730999671692324,
  0.113462997762777, -0.112847998000707, 0.161617065299512,
  0.0417842527227712, 0.0109339973072024, 0.0873866020462818,
  -0.313518196763554, 0.495209512276699, -0.557565321921219,
  0.970467311515782, -0.0355375332851829, 0.118608040240739,
  -0.206810923131812, -0.355569895276308, -0.0697349025274193,
  -0.961253556513966, -0.929149143871644, 0.249854431575179,
  0.893303290452704, -0.364892856721843, 0.0979906699009544,
  -0.27362395883046, 0.145610986528573, -0.067017735101995,
  -0.331651309255641, 0.35877447250923, 0.164991738131823,
  -0.542544977767251, -0.953628463765595, -1.90386582019867,
  0.236119869941792, -0.287518573062719, -0.181517256455921,
  1.55856055254855, 0.516439274402045, -1.17570012741235,
  0.116471889724383, -1.2651273374079, -0.327328496010877,
  0.00559255448856064, 0.0255997544666548, 0.436392616780441,
  -0.428949930298353, 0.676593273818505, 0.376276455095621,
  0.540695863755132, -0.145074339054826, 0.338907653438328,
  0.132996176038587, -0.430794880583753, 0.241514033446405,
  -0.298688862903542, 0.800210327783666, -0.209584763143457,
  -0.0495087375595963, -0.0975630048461466, 0.00861616907747728,
  0.086859241506515, 0.0044587652258629, -0.0418989610640676,
  -0.669755627116209, -0.826831947078139, -0.0635059333821397,
  0.249585367285994, 0.00558291811915919, 0.546377399105633,
  -0.176296245779617, 0.127332693491771, 0.0587819650465473,
  -0.119841084534812, 1.17999885523759, -0.848544719833527,
  -0.0109753488162034, 0.0644354636195647, -0.691412631878793,
  0.209591725650749, -0.0692485220800213, -0.238358294938817,
  0.305282385721245, 0.97756907187131, -1.11872961789879,
  0.741291018625425, -0.989701612162464, 0.376689094817301,
  -0.00766097213051119, 0.277472260392479, 0.167387856294492,
  -0.631111198983839, 0.875305788398969, -0.125744681740375,
  -0.755369600026632, 1.76486571948705, 0.325930962432382,
  0.0562956910371368, 0.0555662077044383, -0.132507060024583,
  0.284224022069574, -0.349205712020249, -1.01829540069731,
  0.0308222476562478, 0.105235902372921, 0.12629983819838,
  -0.296656450451795, -0.038138154763896, -0.194346220970277,
  -0.421838762145911, 0.463454570343692, -0.36577043603591,
  0.118198413692332, -0.394830515755158, 0.54853434910693,
  -0.348705674469222, -0.306360268493902, -0.0910784899023358,
  -0.198656328297743, 0.514035878160728, 0.45802285990493,
  -0.25805561598919, 0.14861454342082, 0.344776392298896,
  0.021005719854877, 0.0757629480750393, 0.0047098998280666,
  -0.112665516455951, 0.245788710802021, 0.0324571326187557,
  0.0386622675204586, 1.35257649155514, 0.231476620786973,
  -0.166498074336848, -0.129383568567935, -0.145938972600868,
  -0.0278240573418748, 0.0189691193837534, 0.00333524117304829,
  -0.0126222032405218, 0.0068937476384311, -0.0800957394144725,
  0.0802332309514961, 0.234983482044546, -0.383199046059846,
  0.568488183545177, 1.0327656507292, -1.60066949181259,
  -0.38851294939742, -0.738765575912372, 1.30901544387702,
  -0.0717045883729113, -0.205454153590326, -0.0400329945205947,
  -0.754366101407317, -0.11117381903109, 0.309196425293675,
  -0.204311204324809, 0.643450194765779, -0.047534937415621,
  0.284764206324933, 0.258458530481182, 0.0763695450944505,
  0.279892985117472, 1.14152294975613, -0.372025159471505,
  0.608449851362017, 1.14053242739383, 0.493735544791118,
  -0.011662775833786, -0.212836717261086, 0.0827880258161556,
  -0.631238375566844, -0.631876956551708, 0.0147663872359829,
  -0.817078337500636, -0.766058670649528, -0.0348401341263962,
  -0.0852322772115565, -0.164083573806344, 0.0994339885082557,
  -0.621020867004594, 0.487970188712165, -0.195651723595036,
  0.112650219107924, -0.397999260964717, 1.2632381384419,
  -0.089145313658172, -0.0894304753369774, -0.456330532886704,
  0.154034402767617, -0.604611018240219, 0.939070657411948,
  -0.0578647759228205, 0.13784813509231, -0.887426903413123,
  0.220521557264538, -0.0390066288882564, 0.151647585889686,
  0.157221931817462, 0.321379792700527, 0.303971545292033,
  -1.03772338014671, 0.840398142012763, -0.804248463669083,
  0.0993124847055766, -0.0970866861509242, -0.0285257580968574,
  -0.69677555801569, -0.0672809080358111, -0.431755464936127,
  -0.667978886605616, -0.446353796943168, -0.925780275264681,
  -0.153811026815025, -0.347162700927055, -0.0239608605912896,
  -0.0889543965573955, -0.383299459538774, -0.361427085293351,
  0.208954601737557, 0.331911050292229, 0.280446033259532,
  0.136378338472505, 0.0799027126080594, 0.0129389493698877,
  0.0915546850949052, 0.640919637794064, 0.902180099578664,
  0.121677335964535, -0.575046400441408, -0.276348748014119,
  -0.0358454337925655, 0.2046150819037, -0.0901090155718139,
  -0.0485379369807913, 0.425079441109613, 0.0564103507735586,
  0.16196035709142, -0.219551206047164, -0.189530710706645,
  0.379168722249477, -0.253733915127216, 0.125267729971722,
  -0.847400555347316, 0.249779915633094, -0.277704621150973,
  0.49889566452289, -0.105366272828763, 1.4705148494632,
  0.0868744135004567, 0.142244947649631, 0.148053688476552,
  -0.217016848207455, 0.120704758269749, 0.293656590609841,
  1.12508281999824, 0.15366377077372, 0.441711173126659,
  0.25236386651259, 0.225297139060153, -0.0655329758120583,
  -0.119705606687929, 0.429789502526318, -0.566117040750032,
  -1.00572114011116, -0.375472688722192, 0.965603592718735,
  0.289125546355131, -0.0826350594404479, 0.155048330571595,
  0.328552448777865, -0.225224089598033, -0.00973988621563427,
  0.133745012285267, 0.0965873542197232, 0.0820952058267112,
  -0.161829068646148, 0.117800537404605, -0.176931866393475,
  0.627271185574049, -0.205471387425923, 0.929893956507948,
  -0.416282873858776, 0.798599305445064, 0.0672596559017571,
  0.198282913549976, -0.140689329355541, 0.12588252211515,
  0.484658475288452, -0.68862958991441, 0.344683687630109,
  -0.526771869394222, -0.057494944225573, 0.412061286109985,
  -0.228341038738954, 0.260342006891256, -0.178939608895562,
  -0.417031038767709, 0.000720461458991698, -0.210164578257806,
  -0.529329039085494, 1.31397966501617, 0.0351118139107122,
  -0.0265560466187338, -0.272619853973099, -0.456670994988454,
  0.108063592029535, -0.267472910891646, -0.101943715961704,
  0.03884378046657, -0.124811772388617, -0.877364047872146,
  0.0991092809119278, -0.246718430818099, -0.0946227085340088,
  -0.373444256654788, 0.592713962908651, 0.565526879863198,
  -0.367098658134207, 0.351545700534717, 0.590290700551054,
  -0.145208898607332, -0.183308884804683, 0.0221216049624343,
  -0.0382244105647031, -0.494770484229957, -0.229943339127264,
  0.120708441123341, 0.163863296152566, -0.460068736680899,
  -0.249432885267174, -0.149851990746015, 0.100924793336167,
  -0.439776516578992, 0.0552312443264442, 0.231113185287227,
  0.684966834410217, -0.272339811774831, -0.841592666619969,
  0.191179879390408, -0.124358543092312, 0.156378032685079,
  0.148799575727893, 0.08396842301226, 0.347241001793077,
  0.670398541705696, -1.47165667133187, -0.0718446780263824,
  0.0110831785689567, -0.399431984907493, 0.121785737369718,
  0.391530064482265, 0.39981676006206, -0.244787697271361,
  0.569943613428441, -1.12193671556171, -0.00695010635251444,
  0.248455332425447, 0.0534789687225097, -0.175376943735574,
  -1.30076811149016, -0.197869035924901, -0.323720078886722,
  0.74914499792668, 0.125906377020262, 0.35796889929944,
  0.169907867421492, 0.0809220583648345, -0.037988877028293,
  -0.168658532939469, -0.101352920099595, -0.38062584220423,
  0.021993748560763, 0.0181267475128731, -0.204956588943909,
  0.041964862028234, 0.24550188304049, -0.0122698241281634,
  0.179452603718771, -1.11720522705365, -0.398975326033384,
  0.269670274708847, 0.35222621410982, 0.19111460099103,
  -0.252731096210632, 0.0741819013779072, 0.0321824592760361,
  -0.159341461464212, -0.733506902511536, -0.269669389922483,
  0.132180207650926, 0.484893497937167, 0.566370124633658,
  -0.0779069897666886, -0.220659791343036, -0.251441657719281,
  -0.124450760306334, 0.151341008759725, 0.0449156430853597,
  -0.258235410860573, 0.358993681942866, 0.286392168205914,
  0.0561136448629831, -0.0759758549610551, 0.205476739241104,
  -0.425025132960902, -0.448068691191524, 0.952333040018811,
  0.583181876092715, 0.664917821091343, -1.07141001929735,
  0.316402727372656, 0.378404681076651, -0.338763714228794,
  0.348903242126211, 0.445012446800056, -0.445302364074697,
  0.242177154341399, 0.307311350525707, -0.258192798290928,
  -0.27672003312879, -0.00795975651102303, -0.164608423448828,
  -0.780141421690648, -0.0598598388563096, -1.20671846251848,
  -0.210613727861141, 0.478503415381108, -0.217498856700077,
  0.220048590951193, -0.209637674490311, -0.276187854583098,
  -0.303180635911122, -0.633017835447315, -0.129796965702467,
  0.681040024031705, 0.51469026010616, -0.330517955522662,
  -0.332014933593799, 0.407338391426003, 0.108231603661128,
  -0.729132144414724, 0.028070282775225, -0.283994621872146,
  0.319885744990133, 0.576544467007221, 0.341191636546231,
  -0.2404223351243, 0.114564852543929, 0.119497271589942,
  -0.598712869200023, -1.04644457258893, -0.492275478152766,
  0.101534590295471, 0.474969383274721, 0.182819441964283,
  -0.117096066154396, -0.0600845663205416, 0.0698050276684972,
  -0.464746720370855, 1.05992655159159, -0.506849453284128,
  -0.258407889638925, 0.597159216249164, -0.251040159303181,
  -0.137422442863663, 0.224587329334157, -0.0434861811163645,
  -0.36648727972605, -0.0696816571483855, 0.369753875445986,
  -1.24995929521305, 0.223334038906147, 0.703238902956571,
  -0.247409886496191, -0.111542996763804, -0.00200854033163777,
  -0.507252118195684, 0.254410899283535, 0.0397871085227668,
  -0.523680209417583, 0.114997549262223, -0.20356261999245,
  0.159329695416569, 0.209432720183252, 0.0207597952564806,
  0.242096644196771, -0.34722986059327, 0.192218801014268,
  0.406101831447595, 0.0476450492823598, -0.946340927072305,
  0.0455547308241934, -0.0395532518160629, 0.0527652915552157,
  -0.138734204835149, 0.149510252081293, -0.282034388079668,
  -0.036215648977248, -0.786993287484684, 0.739843769689148,
  0.0702062400335691, -0.288150937377671, 0.104874922767834,
  -0.155451155894122, 0.169389538118713, -0.139802487353832,
  0.0850893821465697, -0.0421407868933928, -0.00320959265492306,
  0.379290574409844, 0.252312107003208, 0.0958436328184011,
  0.956096306352713, 0.15857917957553, -1.59460393776291,
  -0.768103430482038, 1.60972167432007, 0.257323789791101,
  -0.125879660191345, -0.00806100246015264, 0.310334009256379,
  -0.627139172790466, -0.49113933878432, 0.602899824550157,
  0.0636799955478798, -0.269102037167718, 0.860821561293212,
  -0.285720817048907, 0.100954338601068, -0.198244706012297,
  -0.260160847147215, 0.642411959402278, -0.686476137314227,
  0.870294355632454, 0.499102866039368, 1.25290294343595,
  0.0401973857540271, -0.224939309281113, -0.167331825059847,
  0.336195021038107, 0.504075906382392, 0.210859451415977,
  -0.297078998716589, 0.134012442021256, -0.147159916165614,
  0.192058845745943, 0.109731912251015, -0.101153317235968,
  0.496057951148426, 0.647377128193584, -0.361785291927689,
  0.465826442721069, -0.29782111105142, -0.801780410524583,
  -0.122762325489805, 0.0835967652895686, 0.0306842883101144,
  -0.101623294593458, -0.141308234027055, -0.00984859168712517,
  1.13093688416115, 0.363769375206935, 0.287017625357163,
  -0.12164691393067, 0.0952179448437575, -0.0198600461761554,
  -0.216837161516116, 0.857848341081296, -0.0551447598247526,
  0.0478435182183467, 1.00724822403552, -0.0507932588419517,
  -0.0958526882825772, -0.0825850492733874, 0.0600191838359879,
  -0.423918064674118, 0.980442460061949, -0.252505945079693,
  0.532075366560572, -1.06773717912419, 0.309797673121148,
  0.289632857537965, 0.266360126341266, -0.0763221824804867,
  -0.233910100881588, -0.0641454812587651, -0.18665715708,
  0.267482863485978, 0.721117421163012, -0.460561074753846,
  -0.269349882429433, -0.0452088267878307, -0.00599606172306296,
  -0.240381945991158, 0.0604266494938889, -0.245609070613803,
  -0.467513947442889, 0.0773601638785848, 0.119075022975661,
  0.304869895136032, 0.0397340158500657, -0.274807773549111,
  -0.977607235463285, 0.391438267553967, -0.92437201772607,
  0.485218659819626, -0.150617599140947, -0.0660040102485444,
  -0.128971861417356, -0.102298124682158, 0.221715929456246,
  -0.094601206545487, -0.242704872970128, -0.225565995953185,
  -0.188389677602765, 0.00223485054891892, 0.542190294504877,
  0.154705296350126, -0.10509263946069, 0.332448929027376,
  0.0264585221267943, 0.125288033921623, 0.152401940571733,
  -0.219272422399779, 0.0724531516481246, -0.802255639832044,
  -0.347597469034255, -0.033580815012224, -0.17662338802779,
  -1.0041176426334, 0.37587378803889, -0.474125812198235,
  -0.275147747329801, -0.18494538263267, -0.132986812571721,
  0.105507169120013, 0.0484690298010166, 0.0714879429213614,
  0.0546335243461732, 0.05619242327035, -0.133512927015966,
  0.953029532475567, 1.33647865358866, 0.474781792609853,
  -0.335321824203395, -0.186779201430801, -0.102932062747404,
  -0.927789020287163, -0.851327699536668, -0.636246409128869,
  -0.807270538046092, 0.457808777018289, 0.240436354895732,
  -0.31149989927279, -0.0416306098624421, -0.239061492515207,
  0.225783582215596, 0.060302836463749, -0.279368729776076,
  -0.46440797716751, -0.312260488881195, -0.875472932358936,
  -0.0330204107764939, -0.162749846902038, 0.260119029658435,
  0.147004640450984, -0.0587995982512783, 0.167026965965079,
  -0.0730106305227905, 0.00568973089906798, 0.319038498205732,
  -0.103270532724575, -0.0692147169199323, 0.00552852757710388,
  0.152117458267483, 0.520069001568054, -0.580103265733194,
  -0.166420881962733, 0.515171218007504, 0.0861507127814736,
  -0.224842148605954, 0.112095097092397, 0.131546957996599,
  -0.876773859248005, 0.544584347466835, -0.417827971688385,
  0.362581590074217, -0.526896360250131, 0.767220497264671,
  -0.533621731666685, -0.215069089731718, -0.237303055795645,
  1.02115968180952, 1.3980912866903, -0.598398555235081,
  -0.985540246000373, 1.06410647164351, 0.572379240043525,
  -0.0021596112556583, 0.0349183542936309, -0.0515575903012726,
  0.354967077756763, 0.0715447495028106, 0.371590116783388,
  0.487491527052814, -0.0393808586290617, -0.753067695825824,
  -0.0037761191653331, -0.260945920839552, 0.0162282190191539,
  0.618207658145769, -0.663171035021779, 0.0924276647387517,
  -0.0877321709536261, 0.0761008997276113, -0.0733813913452413,
  -0.238534713955533, 0.117999336780344, 0.0988294076896362,
  -0.00915865077207889, -0.579867115553333, -0.214275202213707,
  -0.39888391772915, 0.314258716816458, 0.161363198132749,
  0.442805919080865, 0.0605206603039656, 0.16265789641071,
  0.570544758495884, -0.702611915237217, -0.591172202468745,
  -1.27112721085449, 0.336654990311977, 0.38166423262562,
  -0.125057565181075, -0.162443237220827, 0.100833088811078,
  -0.2752337450214, -0.380414809972686, 0.422112402472388,
  1.47968139660452, -0.358572736322888, 0.881334207356249,
  -0.0306828632797499, 0.346726157354006, 0.0984324120736902,
  -0.0721034992777305, -0.0984880387196832, -0.691588086951366,
  0.451835047250376, -0.870710290490948, 0.156857821149449,
  -0.109463623005918, 0.00714598040510136, -0.145482831294702,
  -0.0396818514545868, 0.319460198364389, -0.117382329996837,
  0.135871941632839, -0.00737825195149069, 0.974924926811074,
  -0.031715103290114, -0.0431204135765418, -3.0356316487672275,
  -0.00155236562319001, -0.357499640488191, -3.1489187360697060,
  -0.0909185010127125, 0.360084667499076, -3.214425116585007 ;

 cell_spatial = "abc" ;

 cell_angular =
  "alpha",
  "beta ",
  "gamma" ;

 cell_lengths = 31.077, 31.077, 150 ;

 cell_angles = 90, 90, 90 ;
}
